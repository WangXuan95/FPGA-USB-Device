
//--------------------------------------------------------------------------------------------------------
// Module  : fpga_top_usb_disk
// Type    : synthesizable, fpga top
// Standard: Verilog 2001 (IEEE1364-2001)
// Function: example for usb_disk_top
//--------------------------------------------------------------------------------------------------------

module fpga_top_usb_disk (
    // clock
    input  wire        clk50mhz,     // connect to a 50MHz oscillator
    // reset button
    input  wire        button,       // connect to a reset button, 0=reset, 1=release. If you don't have a button, tie this signal to 1.
    // LED
    output wire        led,          // 1: USB connected , 0: USB disconnected
    // USB signals
    output wire        usb_dp_pull,  // connect to USB D+ by an 1.5k resistor
    inout              usb_dp,       // connect to USB D+
    inout              usb_dn,       // connect to USB D-
    // debug output info, only for USB developers, can be ignored for normally use
    output wire        uart_tx       // If you want to see the debug info of USB device core, please connect this UART signal to host-PC (UART format: 115200,8,n,1), otherwise you can ignore this signal.
);




//-------------------------------------------------------------------------------------------------------------------------------------
// The USB controller core needs a 60MHz clock, this PLL module is to convert clk50mhz to clk60mhz
// This PLL module is only available on Altera Cyclone IV E.
// If you use other FPGA families, please use their compatible primitives or IP-cores to generate clk60mhz
//-------------------------------------------------------------------------------------------------------------------------------------
wire [3:0] subwire0;
wire       clk60mhz;
wire       clk_locked;
altpll u_altpll (
    .inclk       ( {1'b0, clk50mhz}     ),
    .clk         ( {subwire0, clk60mhz} ),
    .locked      ( clk_locked           ),
    .activeclock (),    .areset (1'b0),    .clkbad (),    .clkena ({6{1'b1}}),    .clkloss (),    .clkswitch (1'b0),    .configupdate (1'b0),    .enable0 (),    .enable1 (),    .extclk (),    .extclkena ({4{1'b1}}),    .fbin (1'b1),    .fbmimicbidir (),    .fbout (),    .fref (),    .icdrclk (),    .pfdena (1'b1),    .phasecounterselect ({4{1'b1}}),    .phasedone (),    .phasestep (1'b1),    .phaseupdown (1'b1),    .pllena (1'b1),    .scanaclr (1'b0),    .scanclk (1'b0),    .scanclkena (1'b1),    .scandata (1'b0),    .scandataout (),    .scandone (),    .scanread (1'b0),    .scanwrite (1'b0),    .sclkout0 (),    .sclkout1 (),    .vcooverrange (),    .vcounderrange () );
defparam u_altpll.bandwidth_type = "AUTO",    u_altpll.clk0_divide_by = 5,    u_altpll.clk0_duty_cycle = 50,    u_altpll.clk0_multiply_by = 6,    u_altpll.clk0_phase_shift = "0",    u_altpll.compensate_clock = "CLK0",    u_altpll.inclk0_input_frequency = 20000,    u_altpll.intended_device_family = "Cyclone IV E",    u_altpll.lpm_hint = "CBX_MODULE_PREFIX=pll",    u_altpll.lpm_type = "altpll",    u_altpll.operation_mode = "NORMAL",    u_altpll.pll_type = "AUTO",    u_altpll.port_activeclock = "PORT_UNUSED",    u_altpll.port_areset = "PORT_UNUSED",    u_altpll.port_clkbad0 = "PORT_UNUSED",    u_altpll.port_clkbad1 = "PORT_UNUSED",    u_altpll.port_clkloss = "PORT_UNUSED",    u_altpll.port_clkswitch = "PORT_UNUSED",    u_altpll.port_configupdate = "PORT_UNUSED",    u_altpll.port_fbin = "PORT_UNUSED",    u_altpll.port_inclk0 = "PORT_USED",    u_altpll.port_inclk1 = "PORT_UNUSED",    u_altpll.port_locked = "PORT_USED",    u_altpll.port_pfdena = "PORT_UNUSED",    u_altpll.port_phasecounterselect = "PORT_UNUSED",    u_altpll.port_phasedone = "PORT_UNUSED",    u_altpll.port_phasestep = "PORT_UNUSED",    u_altpll.port_phaseupdown = "PORT_UNUSED",    u_altpll.port_pllena = "PORT_UNUSED",    u_altpll.port_scanaclr = "PORT_UNUSED",    u_altpll.port_scanclk = "PORT_UNUSED",    u_altpll.port_scanclkena = "PORT_UNUSED",    u_altpll.port_scandata = "PORT_UNUSED",    u_altpll.port_scandataout = "PORT_UNUSED",    u_altpll.port_scandone = "PORT_UNUSED",    u_altpll.port_scanread = "PORT_UNUSED",    u_altpll.port_scanwrite = "PORT_UNUSED",    u_altpll.port_clk0 = "PORT_USED",    u_altpll.port_clk1 = "PORT_UNUSED",    u_altpll.port_clk2 = "PORT_UNUSED",    u_altpll.port_clk3 = "PORT_UNUSED",    u_altpll.port_clk4 = "PORT_UNUSED",    u_altpll.port_clk5 = "PORT_UNUSED",    u_altpll.port_clkena0 = "PORT_UNUSED",    u_altpll.port_clkena1 = "PORT_UNUSED",    u_altpll.port_clkena2 = "PORT_UNUSED",    u_altpll.port_clkena3 = "PORT_UNUSED",    u_altpll.port_clkena4 = "PORT_UNUSED",    u_altpll.port_clkena5 = "PORT_UNUSED",    u_altpll.port_extclk0 = "PORT_UNUSED",    u_altpll.port_extclk1 = "PORT_UNUSED",    u_altpll.port_extclk2 = "PORT_UNUSED",    u_altpll.port_extclk3 = "PORT_UNUSED",    u_altpll.self_reset_on_loss_lock = "OFF",    u_altpll.width_clock = 5;




//-------------------------------------------------------------------------------------------------------------------------------------
// USB-MSC disk device
//-------------------------------------------------------------------------------------------------------------------------------------

wire [40:0] mem_addr;
wire        mem_wen;
wire [ 7:0] mem_wdata;
reg  [ 7:0] mem_rdata;

usb_disk_top #(
    .BLOCK_COUNT     ( 48                  ),   // block count of the disk, each block has 512 bytes. Here it has 48 blocks = 24kiB
    .DEBUG           ( "FALSE"             )    // If you want to see the debug info of USB device core, set this parameter to "TRUE"
) u_usb_disk (
    .rstn            ( clk_locked & button ),
    .clk             ( clk60mhz            ),
    // USB signals
    .usb_dp_pull     ( usb_dp_pull         ),
    .usb_dp          ( usb_dp              ),
    .usb_dn          ( usb_dn              ),
    // USB reset output
    .usb_rstn        ( led                 ),   // 1: connected , 0: disconnected (when USB cable unplug, or when system reset (rstn=0))
    // disk memory access interface
    .mem_addr        ( mem_addr            ),   // byte address
    .mem_wen         ( mem_wen             ),   // 1:write   0:read
    .mem_wdata       ( mem_wdata           ),   // byte to write
    .mem_rdata       ( mem_rdata           ),   // byte to read
    // debug output info, only for USB developers, can be ignored for normally use
    .debug_en        (                     ),
    .debug_data      (                     ),
    .debug_uart_tx   ( uart_tx             )
);




//-------------------------------------------------------------------------------------------------------------------------------------
// a 24kiB disk memory (implement with BRAM), the initial values contain a simple FAT file-system
//-------------------------------------------------------------------------------------------------------------------------------------
reg [7:0] disk_mem [0:24575];
always @ (posedge clk60mhz) mem_rdata <= disk_mem[mem_addr[14:0]];
always @ (posedge clk60mhz) if(mem_wen)  disk_mem[mem_addr[14:0]] <= mem_wdata;


initial begin
disk_mem[    0] = 0;
disk_mem[    1] = 0;
disk_mem[    2] = 0;
disk_mem[    3] = 0;
disk_mem[    4] = 0;
disk_mem[    5] = 0;
disk_mem[    6] = 0;
disk_mem[    7] = 0;
disk_mem[    8] = 0;
disk_mem[    9] = 0;
disk_mem[   10] = 0;
disk_mem[   11] = 0;
disk_mem[   12] = 0;
disk_mem[   13] = 0;
disk_mem[   14] = 0;
disk_mem[   15] = 0;
disk_mem[   16] = 0;
disk_mem[   17] = 0;
disk_mem[   18] = 0;
disk_mem[   19] = 0;
disk_mem[   20] = 0;
disk_mem[   21] = 0;
disk_mem[   22] = 0;
disk_mem[   23] = 0;
disk_mem[   24] = 0;
disk_mem[   25] = 0;
disk_mem[   26] = 0;
disk_mem[   27] = 0;
disk_mem[   28] = 0;
disk_mem[   29] = 0;
disk_mem[   30] = 0;
disk_mem[   31] = 0;
disk_mem[   32] = 0;
disk_mem[   33] = 0;
disk_mem[   34] = 0;
disk_mem[   35] = 0;
disk_mem[   36] = 0;
disk_mem[   37] = 0;
disk_mem[   38] = 0;
disk_mem[   39] = 0;
disk_mem[   40] = 0;
disk_mem[   41] = 0;
disk_mem[   42] = 0;
disk_mem[   43] = 0;
disk_mem[   44] = 0;
disk_mem[   45] = 0;
disk_mem[   46] = 0;
disk_mem[   47] = 0;
disk_mem[   48] = 0;
disk_mem[   49] = 0;
disk_mem[   50] = 0;
disk_mem[   51] = 0;
disk_mem[   52] = 0;
disk_mem[   53] = 0;
disk_mem[   54] = 0;
disk_mem[   55] = 0;
disk_mem[   56] = 0;
disk_mem[   57] = 0;
disk_mem[   58] = 0;
disk_mem[   59] = 0;
disk_mem[   60] = 0;
disk_mem[   61] = 0;
disk_mem[   62] = 0;
disk_mem[   63] = 0;
disk_mem[   64] = 0;
disk_mem[   65] = 0;
disk_mem[   66] = 0;
disk_mem[   67] = 0;
disk_mem[   68] = 0;
disk_mem[   69] = 0;
disk_mem[   70] = 0;
disk_mem[   71] = 0;
disk_mem[   72] = 0;
disk_mem[   73] = 0;
disk_mem[   74] = 0;
disk_mem[   75] = 0;
disk_mem[   76] = 0;
disk_mem[   77] = 0;
disk_mem[   78] = 0;
disk_mem[   79] = 0;
disk_mem[   80] = 0;
disk_mem[   81] = 0;
disk_mem[   82] = 0;
disk_mem[   83] = 0;
disk_mem[   84] = 0;
disk_mem[   85] = 0;
disk_mem[   86] = 0;
disk_mem[   87] = 0;
disk_mem[   88] = 0;
disk_mem[   89] = 0;
disk_mem[   90] = 0;
disk_mem[   91] = 0;
disk_mem[   92] = 0;
disk_mem[   93] = 0;
disk_mem[   94] = 0;
disk_mem[   95] = 0;
disk_mem[   96] = 0;
disk_mem[   97] = 0;
disk_mem[   98] = 0;
disk_mem[   99] = 0;
disk_mem[  100] = 0;
disk_mem[  101] = 0;
disk_mem[  102] = 0;
disk_mem[  103] = 0;
disk_mem[  104] = 0;
disk_mem[  105] = 0;
disk_mem[  106] = 0;
disk_mem[  107] = 0;
disk_mem[  108] = 0;
disk_mem[  109] = 0;
disk_mem[  110] = 0;
disk_mem[  111] = 0;
disk_mem[  112] = 0;
disk_mem[  113] = 0;
disk_mem[  114] = 0;
disk_mem[  115] = 0;
disk_mem[  116] = 0;
disk_mem[  117] = 0;
disk_mem[  118] = 0;
disk_mem[  119] = 0;
disk_mem[  120] = 0;
disk_mem[  121] = 0;
disk_mem[  122] = 0;
disk_mem[  123] = 0;
disk_mem[  124] = 0;
disk_mem[  125] = 0;
disk_mem[  126] = 0;
disk_mem[  127] = 0;
disk_mem[  128] = 0;
disk_mem[  129] = 0;
disk_mem[  130] = 0;
disk_mem[  131] = 0;
disk_mem[  132] = 0;
disk_mem[  133] = 0;
disk_mem[  134] = 0;
disk_mem[  135] = 0;
disk_mem[  136] = 0;
disk_mem[  137] = 0;
disk_mem[  138] = 0;
disk_mem[  139] = 0;
disk_mem[  140] = 0;
disk_mem[  141] = 0;
disk_mem[  142] = 0;
disk_mem[  143] = 0;
disk_mem[  144] = 0;
disk_mem[  145] = 0;
disk_mem[  146] = 0;
disk_mem[  147] = 0;
disk_mem[  148] = 0;
disk_mem[  149] = 0;
disk_mem[  150] = 0;
disk_mem[  151] = 0;
disk_mem[  152] = 0;
disk_mem[  153] = 0;
disk_mem[  154] = 0;
disk_mem[  155] = 0;
disk_mem[  156] = 0;
disk_mem[  157] = 0;
disk_mem[  158] = 0;
disk_mem[  159] = 0;
disk_mem[  160] = 0;
disk_mem[  161] = 0;
disk_mem[  162] = 0;
disk_mem[  163] = 0;
disk_mem[  164] = 0;
disk_mem[  165] = 0;
disk_mem[  166] = 0;
disk_mem[  167] = 0;
disk_mem[  168] = 0;
disk_mem[  169] = 0;
disk_mem[  170] = 0;
disk_mem[  171] = 0;
disk_mem[  172] = 0;
disk_mem[  173] = 0;
disk_mem[  174] = 0;
disk_mem[  175] = 0;
disk_mem[  176] = 0;
disk_mem[  177] = 0;
disk_mem[  178] = 0;
disk_mem[  179] = 0;
disk_mem[  180] = 0;
disk_mem[  181] = 0;
disk_mem[  182] = 0;
disk_mem[  183] = 0;
disk_mem[  184] = 0;
disk_mem[  185] = 0;
disk_mem[  186] = 0;
disk_mem[  187] = 0;
disk_mem[  188] = 0;
disk_mem[  189] = 0;
disk_mem[  190] = 0;
disk_mem[  191] = 0;
disk_mem[  192] = 0;
disk_mem[  193] = 0;
disk_mem[  194] = 0;
disk_mem[  195] = 0;
disk_mem[  196] = 0;
disk_mem[  197] = 0;
disk_mem[  198] = 0;
disk_mem[  199] = 0;
disk_mem[  200] = 0;
disk_mem[  201] = 0;
disk_mem[  202] = 0;
disk_mem[  203] = 0;
disk_mem[  204] = 0;
disk_mem[  205] = 0;
disk_mem[  206] = 0;
disk_mem[  207] = 0;
disk_mem[  208] = 0;
disk_mem[  209] = 0;
disk_mem[  210] = 0;
disk_mem[  211] = 0;
disk_mem[  212] = 0;
disk_mem[  213] = 0;
disk_mem[  214] = 0;
disk_mem[  215] = 0;
disk_mem[  216] = 0;
disk_mem[  217] = 0;
disk_mem[  218] = 0;
disk_mem[  219] = 0;
disk_mem[  220] = 0;
disk_mem[  221] = 0;
disk_mem[  222] = 0;
disk_mem[  223] = 0;
disk_mem[  224] = 0;
disk_mem[  225] = 0;
disk_mem[  226] = 0;
disk_mem[  227] = 0;
disk_mem[  228] = 0;
disk_mem[  229] = 0;
disk_mem[  230] = 0;
disk_mem[  231] = 0;
disk_mem[  232] = 0;
disk_mem[  233] = 0;
disk_mem[  234] = 0;
disk_mem[  235] = 0;
disk_mem[  236] = 0;
disk_mem[  237] = 0;
disk_mem[  238] = 0;
disk_mem[  239] = 0;
disk_mem[  240] = 0;
disk_mem[  241] = 0;
disk_mem[  242] = 0;
disk_mem[  243] = 0;
disk_mem[  244] = 0;
disk_mem[  245] = 0;
disk_mem[  246] = 0;
disk_mem[  247] = 0;
disk_mem[  248] = 0;
disk_mem[  249] = 0;
disk_mem[  250] = 0;
disk_mem[  251] = 0;
disk_mem[  252] = 0;
disk_mem[  253] = 0;
disk_mem[  254] = 0;
disk_mem[  255] = 0;
disk_mem[  256] = 0;
disk_mem[  257] = 0;
disk_mem[  258] = 0;
disk_mem[  259] = 0;
disk_mem[  260] = 0;
disk_mem[  261] = 0;
disk_mem[  262] = 0;
disk_mem[  263] = 0;
disk_mem[  264] = 0;
disk_mem[  265] = 0;
disk_mem[  266] = 0;
disk_mem[  267] = 0;
disk_mem[  268] = 0;
disk_mem[  269] = 0;
disk_mem[  270] = 0;
disk_mem[  271] = 0;
disk_mem[  272] = 0;
disk_mem[  273] = 0;
disk_mem[  274] = 0;
disk_mem[  275] = 0;
disk_mem[  276] = 0;
disk_mem[  277] = 0;
disk_mem[  278] = 0;
disk_mem[  279] = 0;
disk_mem[  280] = 0;
disk_mem[  281] = 0;
disk_mem[  282] = 0;
disk_mem[  283] = 0;
disk_mem[  284] = 0;
disk_mem[  285] = 0;
disk_mem[  286] = 0;
disk_mem[  287] = 0;
disk_mem[  288] = 0;
disk_mem[  289] = 0;
disk_mem[  290] = 0;
disk_mem[  291] = 0;
disk_mem[  292] = 0;
disk_mem[  293] = 0;
disk_mem[  294] = 0;
disk_mem[  295] = 0;
disk_mem[  296] = 0;
disk_mem[  297] = 0;
disk_mem[  298] = 0;
disk_mem[  299] = 0;
disk_mem[  300] = 0;
disk_mem[  301] = 0;
disk_mem[  302] = 0;
disk_mem[  303] = 0;
disk_mem[  304] = 0;
disk_mem[  305] = 0;
disk_mem[  306] = 0;
disk_mem[  307] = 0;
disk_mem[  308] = 0;
disk_mem[  309] = 0;
disk_mem[  310] = 0;
disk_mem[  311] = 0;
disk_mem[  312] = 0;
disk_mem[  313] = 0;
disk_mem[  314] = 0;
disk_mem[  315] = 0;
disk_mem[  316] = 0;
disk_mem[  317] = 0;
disk_mem[  318] = 0;
disk_mem[  319] = 0;
disk_mem[  320] = 0;
disk_mem[  321] = 0;
disk_mem[  322] = 0;
disk_mem[  323] = 0;
disk_mem[  324] = 0;
disk_mem[  325] = 0;
disk_mem[  326] = 0;
disk_mem[  327] = 0;
disk_mem[  328] = 0;
disk_mem[  329] = 0;
disk_mem[  330] = 0;
disk_mem[  331] = 0;
disk_mem[  332] = 0;
disk_mem[  333] = 0;
disk_mem[  334] = 0;
disk_mem[  335] = 0;
disk_mem[  336] = 0;
disk_mem[  337] = 0;
disk_mem[  338] = 0;
disk_mem[  339] = 0;
disk_mem[  340] = 0;
disk_mem[  341] = 0;
disk_mem[  342] = 0;
disk_mem[  343] = 0;
disk_mem[  344] = 0;
disk_mem[  345] = 0;
disk_mem[  346] = 0;
disk_mem[  347] = 0;
disk_mem[  348] = 0;
disk_mem[  349] = 0;
disk_mem[  350] = 0;
disk_mem[  351] = 0;
disk_mem[  352] = 0;
disk_mem[  353] = 0;
disk_mem[  354] = 0;
disk_mem[  355] = 0;
disk_mem[  356] = 0;
disk_mem[  357] = 0;
disk_mem[  358] = 0;
disk_mem[  359] = 0;
disk_mem[  360] = 0;
disk_mem[  361] = 0;
disk_mem[  362] = 0;
disk_mem[  363] = 0;
disk_mem[  364] = 0;
disk_mem[  365] = 0;
disk_mem[  366] = 0;
disk_mem[  367] = 0;
disk_mem[  368] = 0;
disk_mem[  369] = 0;
disk_mem[  370] = 0;
disk_mem[  371] = 0;
disk_mem[  372] = 0;
disk_mem[  373] = 0;
disk_mem[  374] = 0;
disk_mem[  375] = 0;
disk_mem[  376] = 0;
disk_mem[  377] = 0;
disk_mem[  378] = 0;
disk_mem[  379] = 0;
disk_mem[  380] = 0;
disk_mem[  381] = 0;
disk_mem[  382] = 0;
disk_mem[  383] = 0;
disk_mem[  384] = 0;
disk_mem[  385] = 0;
disk_mem[  386] = 0;
disk_mem[  387] = 0;
disk_mem[  388] = 0;
disk_mem[  389] = 0;
disk_mem[  390] = 0;
disk_mem[  391] = 0;
disk_mem[  392] = 0;
disk_mem[  393] = 0;
disk_mem[  394] = 0;
disk_mem[  395] = 0;
disk_mem[  396] = 0;
disk_mem[  397] = 0;
disk_mem[  398] = 0;
disk_mem[  399] = 0;
disk_mem[  400] = 0;
disk_mem[  401] = 0;
disk_mem[  402] = 0;
disk_mem[  403] = 0;
disk_mem[  404] = 0;
disk_mem[  405] = 0;
disk_mem[  406] = 0;
disk_mem[  407] = 0;
disk_mem[  408] = 0;
disk_mem[  409] = 0;
disk_mem[  410] = 0;
disk_mem[  411] = 0;
disk_mem[  412] = 0;
disk_mem[  413] = 0;
disk_mem[  414] = 0;
disk_mem[  415] = 0;
disk_mem[  416] = 0;
disk_mem[  417] = 0;
disk_mem[  418] = 0;
disk_mem[  419] = 0;
disk_mem[  420] = 0;
disk_mem[  421] = 0;
disk_mem[  422] = 0;
disk_mem[  423] = 0;
disk_mem[  424] = 0;
disk_mem[  425] = 0;
disk_mem[  426] = 0;
disk_mem[  427] = 0;
disk_mem[  428] = 0;
disk_mem[  429] = 0;
disk_mem[  430] = 0;
disk_mem[  431] = 0;
disk_mem[  432] = 0;
disk_mem[  433] = 0;
disk_mem[  434] = 0;
disk_mem[  435] = 0;
disk_mem[  436] = 0;
disk_mem[  437] = 0;
disk_mem[  438] = 0;
disk_mem[  439] = 0;
disk_mem[  440] = 'hB3;
disk_mem[  441] = 'h25;
disk_mem[  442] = 'hB9;
disk_mem[  443] = 'h2A;
disk_mem[  444] = 0;
disk_mem[  445] = 0;
disk_mem[  446] = 0;
disk_mem[  447] = 0;
disk_mem[  448] = 'h02;
disk_mem[  449] = 0;
disk_mem[  450] = 'h0E;
disk_mem[  451] = 0;
disk_mem[  452] = 'h30;
disk_mem[  453] = 0;
disk_mem[  454] = 'h01;
disk_mem[  455] = 0;
disk_mem[  456] = 0;
disk_mem[  457] = 0;
disk_mem[  458] = 'h2F;
disk_mem[  459] = 0;
disk_mem[  460] = 0;
disk_mem[  461] = 0;
disk_mem[  462] = 0;
disk_mem[  463] = 0;
disk_mem[  464] = 0;
disk_mem[  465] = 0;
disk_mem[  466] = 0;
disk_mem[  467] = 0;
disk_mem[  468] = 0;
disk_mem[  469] = 0;
disk_mem[  470] = 0;
disk_mem[  471] = 0;
disk_mem[  472] = 0;
disk_mem[  473] = 0;
disk_mem[  474] = 0;
disk_mem[  475] = 0;
disk_mem[  476] = 0;
disk_mem[  477] = 0;
disk_mem[  478] = 0;
disk_mem[  479] = 0;
disk_mem[  480] = 0;
disk_mem[  481] = 0;
disk_mem[  482] = 0;
disk_mem[  483] = 0;
disk_mem[  484] = 0;
disk_mem[  485] = 0;
disk_mem[  486] = 0;
disk_mem[  487] = 0;
disk_mem[  488] = 0;
disk_mem[  489] = 0;
disk_mem[  490] = 0;
disk_mem[  491] = 0;
disk_mem[  492] = 0;
disk_mem[  493] = 0;
disk_mem[  494] = 0;
disk_mem[  495] = 0;
disk_mem[  496] = 0;
disk_mem[  497] = 0;
disk_mem[  498] = 0;
disk_mem[  499] = 0;
disk_mem[  500] = 0;
disk_mem[  501] = 0;
disk_mem[  502] = 0;
disk_mem[  503] = 0;
disk_mem[  504] = 0;
disk_mem[  505] = 0;
disk_mem[  506] = 0;
disk_mem[  507] = 0;
disk_mem[  508] = 0;
disk_mem[  509] = 0;
disk_mem[  510] = 'h55;
disk_mem[  511] = 'hAA;
disk_mem[  512] = 'hEB;
disk_mem[  513] = 'h3C;
disk_mem[  514] = 'h90;
disk_mem[  515] = 'h4D;
disk_mem[  516] = 'h53;
disk_mem[  517] = 'h44;
disk_mem[  518] = 'h4F;
disk_mem[  519] = 'h53;
disk_mem[  520] = 'h35;
disk_mem[  521] = 'h2E;
disk_mem[  522] = 'h30;
disk_mem[  523] = 0;
disk_mem[  524] = 'h02;
disk_mem[  525] = 'h01;
disk_mem[  526] = 'h06;
disk_mem[  527] = 0;
disk_mem[  528] = 'h02;
disk_mem[  529] = 0;
disk_mem[  530] = 'h02;
disk_mem[  531] = 'h2F;
disk_mem[  532] = 0;
disk_mem[  533] = 'hF8;
disk_mem[  534] = 'h01;
disk_mem[  535] = 0;
disk_mem[  536] = 'h3F;
disk_mem[  537] = 0;
disk_mem[  538] = 'hFF;
disk_mem[  539] = 0;
disk_mem[  540] = 'h01;
disk_mem[  541] = 0;
disk_mem[  542] = 0;
disk_mem[  543] = 0;
disk_mem[  544] = 0;
disk_mem[  545] = 0;
disk_mem[  546] = 0;
disk_mem[  547] = 0;
disk_mem[  548] = 'h80;
disk_mem[  549] = 0;
disk_mem[  550] = 'h29;
disk_mem[  551] = 'h81;
disk_mem[  552] = 'h88;
disk_mem[  553] = 'hC5;
disk_mem[  554] = 'h9E;
disk_mem[  555] = 'h4E;
disk_mem[  556] = 'h4F;
disk_mem[  557] = 'h20;
disk_mem[  558] = 'h4E;
disk_mem[  559] = 'h41;
disk_mem[  560] = 'h4D;
disk_mem[  561] = 'h45;
disk_mem[  562] = 'h20;
disk_mem[  563] = 'h20;
disk_mem[  564] = 'h20;
disk_mem[  565] = 'h20;
disk_mem[  566] = 'h46;
disk_mem[  567] = 'h41;
disk_mem[  568] = 'h54;
disk_mem[  569] = 'h31;
disk_mem[  570] = 'h32;
disk_mem[  571] = 'h20;
disk_mem[  572] = 'h20;
disk_mem[  573] = 'h20;
disk_mem[  574] = 'h33;
disk_mem[  575] = 'hC9;
disk_mem[  576] = 'h8E;
disk_mem[  577] = 'hD1;
disk_mem[  578] = 'hBC;
disk_mem[  579] = 'hF0;
disk_mem[  580] = 'h7B;
disk_mem[  581] = 'h8E;
disk_mem[  582] = 'hD9;
disk_mem[  583] = 'hB8;
disk_mem[  584] = 0;
disk_mem[  585] = 'h20;
disk_mem[  586] = 'h8E;
disk_mem[  587] = 'hC0;
disk_mem[  588] = 'hFC;
disk_mem[  589] = 'hBD;
disk_mem[  590] = 0;
disk_mem[  591] = 'h7C;
disk_mem[  592] = 'h38;
disk_mem[  593] = 'h4E;
disk_mem[  594] = 'h24;
disk_mem[  595] = 'h7D;
disk_mem[  596] = 'h24;
disk_mem[  597] = 'h8B;
disk_mem[  598] = 'hC1;
disk_mem[  599] = 'h99;
disk_mem[  600] = 'hE8;
disk_mem[  601] = 'h3C;
disk_mem[  602] = 'h01;
disk_mem[  603] = 'h72;
disk_mem[  604] = 'h1C;
disk_mem[  605] = 'h83;
disk_mem[  606] = 'hEB;
disk_mem[  607] = 'h3A;
disk_mem[  608] = 'h66;
disk_mem[  609] = 'hA1;
disk_mem[  610] = 'h1C;
disk_mem[  611] = 'h7C;
disk_mem[  612] = 'h26;
disk_mem[  613] = 'h66;
disk_mem[  614] = 'h3B;
disk_mem[  615] = 'h07;
disk_mem[  616] = 'h26;
disk_mem[  617] = 'h8A;
disk_mem[  618] = 'h57;
disk_mem[  619] = 'hFC;
disk_mem[  620] = 'h75;
disk_mem[  621] = 'h06;
disk_mem[  622] = 'h80;
disk_mem[  623] = 'hCA;
disk_mem[  624] = 'h02;
disk_mem[  625] = 'h88;
disk_mem[  626] = 'h56;
disk_mem[  627] = 'h02;
disk_mem[  628] = 'h80;
disk_mem[  629] = 'hC3;
disk_mem[  630] = 'h10;
disk_mem[  631] = 'h73;
disk_mem[  632] = 'hEB;
disk_mem[  633] = 'h33;
disk_mem[  634] = 'hC9;
disk_mem[  635] = 'h8A;
disk_mem[  636] = 'h46;
disk_mem[  637] = 'h10;
disk_mem[  638] = 'h98;
disk_mem[  639] = 'hF7;
disk_mem[  640] = 'h66;
disk_mem[  641] = 'h16;
disk_mem[  642] = 'h03;
disk_mem[  643] = 'h46;
disk_mem[  644] = 'h1C;
disk_mem[  645] = 'h13;
disk_mem[  646] = 'h56;
disk_mem[  647] = 'h1E;
disk_mem[  648] = 'h03;
disk_mem[  649] = 'h46;
disk_mem[  650] = 'h0E;
disk_mem[  651] = 'h13;
disk_mem[  652] = 'hD1;
disk_mem[  653] = 'h8B;
disk_mem[  654] = 'h76;
disk_mem[  655] = 'h11;
disk_mem[  656] = 'h60;
disk_mem[  657] = 'h89;
disk_mem[  658] = 'h46;
disk_mem[  659] = 'hFC;
disk_mem[  660] = 'h89;
disk_mem[  661] = 'h56;
disk_mem[  662] = 'hFE;
disk_mem[  663] = 'hB8;
disk_mem[  664] = 'h20;
disk_mem[  665] = 0;
disk_mem[  666] = 'hF7;
disk_mem[  667] = 'hE6;
disk_mem[  668] = 'h8B;
disk_mem[  669] = 'h5E;
disk_mem[  670] = 'h0B;
disk_mem[  671] = 'h03;
disk_mem[  672] = 'hC3;
disk_mem[  673] = 'h48;
disk_mem[  674] = 'hF7;
disk_mem[  675] = 'hF3;
disk_mem[  676] = 'h01;
disk_mem[  677] = 'h46;
disk_mem[  678] = 'hFC;
disk_mem[  679] = 'h11;
disk_mem[  680] = 'h4E;
disk_mem[  681] = 'hFE;
disk_mem[  682] = 'h61;
disk_mem[  683] = 'hBF;
disk_mem[  684] = 0;
disk_mem[  685] = 0;
disk_mem[  686] = 'hE8;
disk_mem[  687] = 'hE6;
disk_mem[  688] = 0;
disk_mem[  689] = 'h72;
disk_mem[  690] = 'h39;
disk_mem[  691] = 'h26;
disk_mem[  692] = 'h38;
disk_mem[  693] = 'h2D;
disk_mem[  694] = 'h74;
disk_mem[  695] = 'h17;
disk_mem[  696] = 'h60;
disk_mem[  697] = 'hB1;
disk_mem[  698] = 'h0B;
disk_mem[  699] = 'hBE;
disk_mem[  700] = 'hA1;
disk_mem[  701] = 'h7D;
disk_mem[  702] = 'hF3;
disk_mem[  703] = 'hA6;
disk_mem[  704] = 'h61;
disk_mem[  705] = 'h74;
disk_mem[  706] = 'h32;
disk_mem[  707] = 'h4E;
disk_mem[  708] = 'h74;
disk_mem[  709] = 'h09;
disk_mem[  710] = 'h83;
disk_mem[  711] = 'hC7;
disk_mem[  712] = 'h20;
disk_mem[  713] = 'h3B;
disk_mem[  714] = 'hFB;
disk_mem[  715] = 'h72;
disk_mem[  716] = 'hE6;
disk_mem[  717] = 'hEB;
disk_mem[  718] = 'hDC;
disk_mem[  719] = 'hA0;
disk_mem[  720] = 'hFB;
disk_mem[  721] = 'h7D;
disk_mem[  722] = 'hB4;
disk_mem[  723] = 'h7D;
disk_mem[  724] = 'h8B;
disk_mem[  725] = 'hF0;
disk_mem[  726] = 'hAC;
disk_mem[  727] = 'h98;
disk_mem[  728] = 'h40;
disk_mem[  729] = 'h74;
disk_mem[  730] = 'h0C;
disk_mem[  731] = 'h48;
disk_mem[  732] = 'h74;
disk_mem[  733] = 'h13;
disk_mem[  734] = 'hB4;
disk_mem[  735] = 'h0E;
disk_mem[  736] = 'hBB;
disk_mem[  737] = 'h07;
disk_mem[  738] = 0;
disk_mem[  739] = 'hCD;
disk_mem[  740] = 'h10;
disk_mem[  741] = 'hEB;
disk_mem[  742] = 'hEF;
disk_mem[  743] = 'hA0;
disk_mem[  744] = 'hFD;
disk_mem[  745] = 'h7D;
disk_mem[  746] = 'hEB;
disk_mem[  747] = 'hE6;
disk_mem[  748] = 'hA0;
disk_mem[  749] = 'hFC;
disk_mem[  750] = 'h7D;
disk_mem[  751] = 'hEB;
disk_mem[  752] = 'hE1;
disk_mem[  753] = 'hCD;
disk_mem[  754] = 'h16;
disk_mem[  755] = 'hCD;
disk_mem[  756] = 'h19;
disk_mem[  757] = 'h26;
disk_mem[  758] = 'h8B;
disk_mem[  759] = 'h55;
disk_mem[  760] = 'h1A;
disk_mem[  761] = 'h52;
disk_mem[  762] = 'hB0;
disk_mem[  763] = 'h01;
disk_mem[  764] = 'hBB;
disk_mem[  765] = 0;
disk_mem[  766] = 0;
disk_mem[  767] = 'hE8;
disk_mem[  768] = 'h3B;
disk_mem[  769] = 0;
disk_mem[  770] = 'h72;
disk_mem[  771] = 'hE8;
disk_mem[  772] = 'h5B;
disk_mem[  773] = 'h8A;
disk_mem[  774] = 'h56;
disk_mem[  775] = 'h24;
disk_mem[  776] = 'hBE;
disk_mem[  777] = 'h0B;
disk_mem[  778] = 'h7C;
disk_mem[  779] = 'h8B;
disk_mem[  780] = 'hFC;
disk_mem[  781] = 'hC7;
disk_mem[  782] = 'h46;
disk_mem[  783] = 'hF0;
disk_mem[  784] = 'h3D;
disk_mem[  785] = 'h7D;
disk_mem[  786] = 'hC7;
disk_mem[  787] = 'h46;
disk_mem[  788] = 'hF4;
disk_mem[  789] = 'h29;
disk_mem[  790] = 'h7D;
disk_mem[  791] = 'h8C;
disk_mem[  792] = 'hD9;
disk_mem[  793] = 'h89;
disk_mem[  794] = 'h4E;
disk_mem[  795] = 'hF2;
disk_mem[  796] = 'h89;
disk_mem[  797] = 'h4E;
disk_mem[  798] = 'hF6;
disk_mem[  799] = 'hC6;
disk_mem[  800] = 'h06;
disk_mem[  801] = 'h96;
disk_mem[  802] = 'h7D;
disk_mem[  803] = 'hCB;
disk_mem[  804] = 'hEA;
disk_mem[  805] = 'h03;
disk_mem[  806] = 0;
disk_mem[  807] = 0;
disk_mem[  808] = 'h20;
disk_mem[  809] = 'h0F;
disk_mem[  810] = 'hB6;
disk_mem[  811] = 'hC8;
disk_mem[  812] = 'h66;
disk_mem[  813] = 'h8B;
disk_mem[  814] = 'h46;
disk_mem[  815] = 'hF8;
disk_mem[  816] = 'h66;
disk_mem[  817] = 'h03;
disk_mem[  818] = 'h46;
disk_mem[  819] = 'h1C;
disk_mem[  820] = 'h66;
disk_mem[  821] = 'h8B;
disk_mem[  822] = 'hD0;
disk_mem[  823] = 'h66;
disk_mem[  824] = 'hC1;
disk_mem[  825] = 'hEA;
disk_mem[  826] = 'h10;
disk_mem[  827] = 'hEB;
disk_mem[  828] = 'h5E;
disk_mem[  829] = 'h0F;
disk_mem[  830] = 'hB6;
disk_mem[  831] = 'hC8;
disk_mem[  832] = 'h4A;
disk_mem[  833] = 'h4A;
disk_mem[  834] = 'h8A;
disk_mem[  835] = 'h46;
disk_mem[  836] = 'h0D;
disk_mem[  837] = 'h32;
disk_mem[  838] = 'hE4;
disk_mem[  839] = 'hF7;
disk_mem[  840] = 'hE2;
disk_mem[  841] = 'h03;
disk_mem[  842] = 'h46;
disk_mem[  843] = 'hFC;
disk_mem[  844] = 'h13;
disk_mem[  845] = 'h56;
disk_mem[  846] = 'hFE;
disk_mem[  847] = 'hEB;
disk_mem[  848] = 'h4A;
disk_mem[  849] = 'h52;
disk_mem[  850] = 'h50;
disk_mem[  851] = 'h06;
disk_mem[  852] = 'h53;
disk_mem[  853] = 'h6A;
disk_mem[  854] = 'h01;
disk_mem[  855] = 'h6A;
disk_mem[  856] = 'h10;
disk_mem[  857] = 'h91;
disk_mem[  858] = 'h8B;
disk_mem[  859] = 'h46;
disk_mem[  860] = 'h18;
disk_mem[  861] = 'h96;
disk_mem[  862] = 'h92;
disk_mem[  863] = 'h33;
disk_mem[  864] = 'hD2;
disk_mem[  865] = 'hF7;
disk_mem[  866] = 'hF6;
disk_mem[  867] = 'h91;
disk_mem[  868] = 'hF7;
disk_mem[  869] = 'hF6;
disk_mem[  870] = 'h42;
disk_mem[  871] = 'h87;
disk_mem[  872] = 'hCA;
disk_mem[  873] = 'hF7;
disk_mem[  874] = 'h76;
disk_mem[  875] = 'h1A;
disk_mem[  876] = 'h8A;
disk_mem[  877] = 'hF2;
disk_mem[  878] = 'h8A;
disk_mem[  879] = 'hE8;
disk_mem[  880] = 'hC0;
disk_mem[  881] = 'hCC;
disk_mem[  882] = 'h02;
disk_mem[  883] = 'h0A;
disk_mem[  884] = 'hCC;
disk_mem[  885] = 'hB8;
disk_mem[  886] = 'h01;
disk_mem[  887] = 'h02;
disk_mem[  888] = 'h80;
disk_mem[  889] = 'h7E;
disk_mem[  890] = 'h02;
disk_mem[  891] = 'h0E;
disk_mem[  892] = 'h75;
disk_mem[  893] = 'h04;
disk_mem[  894] = 'hB4;
disk_mem[  895] = 'h42;
disk_mem[  896] = 'h8B;
disk_mem[  897] = 'hF4;
disk_mem[  898] = 'h8A;
disk_mem[  899] = 'h56;
disk_mem[  900] = 'h24;
disk_mem[  901] = 'hCD;
disk_mem[  902] = 'h13;
disk_mem[  903] = 'h61;
disk_mem[  904] = 'h61;
disk_mem[  905] = 'h72;
disk_mem[  906] = 'h0B;
disk_mem[  907] = 'h40;
disk_mem[  908] = 'h75;
disk_mem[  909] = 'h01;
disk_mem[  910] = 'h42;
disk_mem[  911] = 'h03;
disk_mem[  912] = 'h5E;
disk_mem[  913] = 'h0B;
disk_mem[  914] = 'h49;
disk_mem[  915] = 'h75;
disk_mem[  916] = 'h06;
disk_mem[  917] = 'hF8;
disk_mem[  918] = 'hC3;
disk_mem[  919] = 'h41;
disk_mem[  920] = 'hBB;
disk_mem[  921] = 0;
disk_mem[  922] = 0;
disk_mem[  923] = 'h60;
disk_mem[  924] = 'h66;
disk_mem[  925] = 'h6A;
disk_mem[  926] = 0;
disk_mem[  927] = 'hEB;
disk_mem[  928] = 'hB0;
disk_mem[  929] = 'h42;
disk_mem[  930] = 'h4F;
disk_mem[  931] = 'h4F;
disk_mem[  932] = 'h54;
disk_mem[  933] = 'h4D;
disk_mem[  934] = 'h47;
disk_mem[  935] = 'h52;
disk_mem[  936] = 'h20;
disk_mem[  937] = 'h20;
disk_mem[  938] = 'h20;
disk_mem[  939] = 'h20;
disk_mem[  940] = 'h0D;
disk_mem[  941] = 'h0A;
disk_mem[  942] = 'h52;
disk_mem[  943] = 'h65;
disk_mem[  944] = 'h6D;
disk_mem[  945] = 'h6F;
disk_mem[  946] = 'h76;
disk_mem[  947] = 'h65;
disk_mem[  948] = 'h20;
disk_mem[  949] = 'h64;
disk_mem[  950] = 'h69;
disk_mem[  951] = 'h73;
disk_mem[  952] = 'h6B;
disk_mem[  953] = 'h73;
disk_mem[  954] = 'h20;
disk_mem[  955] = 'h6F;
disk_mem[  956] = 'h72;
disk_mem[  957] = 'h20;
disk_mem[  958] = 'h6F;
disk_mem[  959] = 'h74;
disk_mem[  960] = 'h68;
disk_mem[  961] = 'h65;
disk_mem[  962] = 'h72;
disk_mem[  963] = 'h20;
disk_mem[  964] = 'h6D;
disk_mem[  965] = 'h65;
disk_mem[  966] = 'h64;
disk_mem[  967] = 'h69;
disk_mem[  968] = 'h61;
disk_mem[  969] = 'h2E;
disk_mem[  970] = 'hFF;
disk_mem[  971] = 'h0D;
disk_mem[  972] = 'h0A;
disk_mem[  973] = 'h44;
disk_mem[  974] = 'h69;
disk_mem[  975] = 'h73;
disk_mem[  976] = 'h6B;
disk_mem[  977] = 'h20;
disk_mem[  978] = 'h65;
disk_mem[  979] = 'h72;
disk_mem[  980] = 'h72;
disk_mem[  981] = 'h6F;
disk_mem[  982] = 'h72;
disk_mem[  983] = 'hFF;
disk_mem[  984] = 'h0D;
disk_mem[  985] = 'h0A;
disk_mem[  986] = 'h50;
disk_mem[  987] = 'h72;
disk_mem[  988] = 'h65;
disk_mem[  989] = 'h73;
disk_mem[  990] = 'h73;
disk_mem[  991] = 'h20;
disk_mem[  992] = 'h61;
disk_mem[  993] = 'h6E;
disk_mem[  994] = 'h79;
disk_mem[  995] = 'h20;
disk_mem[  996] = 'h6B;
disk_mem[  997] = 'h65;
disk_mem[  998] = 'h79;
disk_mem[  999] = 'h20;
disk_mem[ 1000] = 'h74;
disk_mem[ 1001] = 'h6F;
disk_mem[ 1002] = 'h20;
disk_mem[ 1003] = 'h72;
disk_mem[ 1004] = 'h65;
disk_mem[ 1005] = 'h73;
disk_mem[ 1006] = 'h74;
disk_mem[ 1007] = 'h61;
disk_mem[ 1008] = 'h72;
disk_mem[ 1009] = 'h74;
disk_mem[ 1010] = 'h0D;
disk_mem[ 1011] = 'h0A;
disk_mem[ 1012] = 0;
disk_mem[ 1013] = 0;
disk_mem[ 1014] = 0;
disk_mem[ 1015] = 0;
disk_mem[ 1016] = 0;
disk_mem[ 1017] = 0;
disk_mem[ 1018] = 0;
disk_mem[ 1019] = 'hAC;
disk_mem[ 1020] = 'hCB;
disk_mem[ 1021] = 'hD8;
disk_mem[ 1022] = 'h55;
disk_mem[ 1023] = 'hAA;
disk_mem[ 1024] = 0;
disk_mem[ 1025] = 0;
disk_mem[ 1026] = 0;
disk_mem[ 1027] = 0;
disk_mem[ 1028] = 0;
disk_mem[ 1029] = 0;
disk_mem[ 1030] = 0;
disk_mem[ 1031] = 0;
disk_mem[ 1032] = 0;
disk_mem[ 1033] = 0;
disk_mem[ 1034] = 0;
disk_mem[ 1035] = 0;
disk_mem[ 1036] = 0;
disk_mem[ 1037] = 0;
disk_mem[ 1038] = 0;
disk_mem[ 1039] = 0;
disk_mem[ 1040] = 0;
disk_mem[ 1041] = 0;
disk_mem[ 1042] = 0;
disk_mem[ 1043] = 0;
disk_mem[ 1044] = 0;
disk_mem[ 1045] = 0;
disk_mem[ 1046] = 0;
disk_mem[ 1047] = 0;
disk_mem[ 1048] = 0;
disk_mem[ 1049] = 0;
disk_mem[ 1050] = 0;
disk_mem[ 1051] = 0;
disk_mem[ 1052] = 0;
disk_mem[ 1053] = 0;
disk_mem[ 1054] = 0;
disk_mem[ 1055] = 0;
disk_mem[ 1056] = 0;
disk_mem[ 1057] = 0;
disk_mem[ 1058] = 0;
disk_mem[ 1059] = 0;
disk_mem[ 1060] = 0;
disk_mem[ 1061] = 0;
disk_mem[ 1062] = 0;
disk_mem[ 1063] = 0;
disk_mem[ 1064] = 0;
disk_mem[ 1065] = 0;
disk_mem[ 1066] = 0;
disk_mem[ 1067] = 0;
disk_mem[ 1068] = 0;
disk_mem[ 1069] = 0;
disk_mem[ 1070] = 0;
disk_mem[ 1071] = 0;
disk_mem[ 1072] = 0;
disk_mem[ 1073] = 0;
disk_mem[ 1074] = 0;
disk_mem[ 1075] = 0;
disk_mem[ 1076] = 0;
disk_mem[ 1077] = 0;
disk_mem[ 1078] = 0;
disk_mem[ 1079] = 0;
disk_mem[ 1080] = 0;
disk_mem[ 1081] = 0;
disk_mem[ 1082] = 0;
disk_mem[ 1083] = 0;
disk_mem[ 1084] = 0;
disk_mem[ 1085] = 0;
disk_mem[ 1086] = 0;
disk_mem[ 1087] = 0;
disk_mem[ 1088] = 0;
disk_mem[ 1089] = 0;
disk_mem[ 1090] = 0;
disk_mem[ 1091] = 0;
disk_mem[ 1092] = 0;
disk_mem[ 1093] = 0;
disk_mem[ 1094] = 0;
disk_mem[ 1095] = 0;
disk_mem[ 1096] = 0;
disk_mem[ 1097] = 0;
disk_mem[ 1098] = 0;
disk_mem[ 1099] = 0;
disk_mem[ 1100] = 0;
disk_mem[ 1101] = 0;
disk_mem[ 1102] = 0;
disk_mem[ 1103] = 0;
disk_mem[ 1104] = 0;
disk_mem[ 1105] = 0;
disk_mem[ 1106] = 0;
disk_mem[ 1107] = 0;
disk_mem[ 1108] = 0;
disk_mem[ 1109] = 0;
disk_mem[ 1110] = 0;
disk_mem[ 1111] = 0;
disk_mem[ 1112] = 0;
disk_mem[ 1113] = 0;
disk_mem[ 1114] = 0;
disk_mem[ 1115] = 0;
disk_mem[ 1116] = 0;
disk_mem[ 1117] = 0;
disk_mem[ 1118] = 0;
disk_mem[ 1119] = 0;
disk_mem[ 1120] = 0;
disk_mem[ 1121] = 0;
disk_mem[ 1122] = 0;
disk_mem[ 1123] = 0;
disk_mem[ 1124] = 0;
disk_mem[ 1125] = 0;
disk_mem[ 1126] = 0;
disk_mem[ 1127] = 0;
disk_mem[ 1128] = 0;
disk_mem[ 1129] = 0;
disk_mem[ 1130] = 0;
disk_mem[ 1131] = 0;
disk_mem[ 1132] = 0;
disk_mem[ 1133] = 0;
disk_mem[ 1134] = 0;
disk_mem[ 1135] = 0;
disk_mem[ 1136] = 0;
disk_mem[ 1137] = 0;
disk_mem[ 1138] = 0;
disk_mem[ 1139] = 0;
disk_mem[ 1140] = 0;
disk_mem[ 1141] = 0;
disk_mem[ 1142] = 0;
disk_mem[ 1143] = 0;
disk_mem[ 1144] = 0;
disk_mem[ 1145] = 0;
disk_mem[ 1146] = 0;
disk_mem[ 1147] = 0;
disk_mem[ 1148] = 0;
disk_mem[ 1149] = 0;
disk_mem[ 1150] = 0;
disk_mem[ 1151] = 0;
disk_mem[ 1152] = 0;
disk_mem[ 1153] = 0;
disk_mem[ 1154] = 0;
disk_mem[ 1155] = 0;
disk_mem[ 1156] = 0;
disk_mem[ 1157] = 0;
disk_mem[ 1158] = 0;
disk_mem[ 1159] = 0;
disk_mem[ 1160] = 0;
disk_mem[ 1161] = 0;
disk_mem[ 1162] = 0;
disk_mem[ 1163] = 0;
disk_mem[ 1164] = 0;
disk_mem[ 1165] = 0;
disk_mem[ 1166] = 0;
disk_mem[ 1167] = 0;
disk_mem[ 1168] = 0;
disk_mem[ 1169] = 0;
disk_mem[ 1170] = 0;
disk_mem[ 1171] = 0;
disk_mem[ 1172] = 0;
disk_mem[ 1173] = 0;
disk_mem[ 1174] = 0;
disk_mem[ 1175] = 0;
disk_mem[ 1176] = 0;
disk_mem[ 1177] = 0;
disk_mem[ 1178] = 0;
disk_mem[ 1179] = 0;
disk_mem[ 1180] = 0;
disk_mem[ 1181] = 0;
disk_mem[ 1182] = 0;
disk_mem[ 1183] = 0;
disk_mem[ 1184] = 0;
disk_mem[ 1185] = 0;
disk_mem[ 1186] = 0;
disk_mem[ 1187] = 0;
disk_mem[ 1188] = 0;
disk_mem[ 1189] = 0;
disk_mem[ 1190] = 0;
disk_mem[ 1191] = 0;
disk_mem[ 1192] = 0;
disk_mem[ 1193] = 0;
disk_mem[ 1194] = 0;
disk_mem[ 1195] = 0;
disk_mem[ 1196] = 0;
disk_mem[ 1197] = 0;
disk_mem[ 1198] = 0;
disk_mem[ 1199] = 0;
disk_mem[ 1200] = 0;
disk_mem[ 1201] = 0;
disk_mem[ 1202] = 0;
disk_mem[ 1203] = 0;
disk_mem[ 1204] = 0;
disk_mem[ 1205] = 0;
disk_mem[ 1206] = 0;
disk_mem[ 1207] = 0;
disk_mem[ 1208] = 0;
disk_mem[ 1209] = 0;
disk_mem[ 1210] = 0;
disk_mem[ 1211] = 0;
disk_mem[ 1212] = 0;
disk_mem[ 1213] = 0;
disk_mem[ 1214] = 0;
disk_mem[ 1215] = 0;
disk_mem[ 1216] = 0;
disk_mem[ 1217] = 0;
disk_mem[ 1218] = 0;
disk_mem[ 1219] = 0;
disk_mem[ 1220] = 0;
disk_mem[ 1221] = 0;
disk_mem[ 1222] = 0;
disk_mem[ 1223] = 0;
disk_mem[ 1224] = 0;
disk_mem[ 1225] = 0;
disk_mem[ 1226] = 0;
disk_mem[ 1227] = 0;
disk_mem[ 1228] = 0;
disk_mem[ 1229] = 0;
disk_mem[ 1230] = 0;
disk_mem[ 1231] = 0;
disk_mem[ 1232] = 0;
disk_mem[ 1233] = 0;
disk_mem[ 1234] = 0;
disk_mem[ 1235] = 0;
disk_mem[ 1236] = 0;
disk_mem[ 1237] = 0;
disk_mem[ 1238] = 0;
disk_mem[ 1239] = 0;
disk_mem[ 1240] = 0;
disk_mem[ 1241] = 0;
disk_mem[ 1242] = 0;
disk_mem[ 1243] = 0;
disk_mem[ 1244] = 0;
disk_mem[ 1245] = 0;
disk_mem[ 1246] = 0;
disk_mem[ 1247] = 0;
disk_mem[ 1248] = 0;
disk_mem[ 1249] = 0;
disk_mem[ 1250] = 0;
disk_mem[ 1251] = 0;
disk_mem[ 1252] = 0;
disk_mem[ 1253] = 0;
disk_mem[ 1254] = 0;
disk_mem[ 1255] = 0;
disk_mem[ 1256] = 0;
disk_mem[ 1257] = 0;
disk_mem[ 1258] = 0;
disk_mem[ 1259] = 0;
disk_mem[ 1260] = 0;
disk_mem[ 1261] = 0;
disk_mem[ 1262] = 0;
disk_mem[ 1263] = 0;
disk_mem[ 1264] = 0;
disk_mem[ 1265] = 0;
disk_mem[ 1266] = 0;
disk_mem[ 1267] = 0;
disk_mem[ 1268] = 0;
disk_mem[ 1269] = 0;
disk_mem[ 1270] = 0;
disk_mem[ 1271] = 0;
disk_mem[ 1272] = 0;
disk_mem[ 1273] = 0;
disk_mem[ 1274] = 0;
disk_mem[ 1275] = 0;
disk_mem[ 1276] = 0;
disk_mem[ 1277] = 0;
disk_mem[ 1278] = 0;
disk_mem[ 1279] = 0;
disk_mem[ 1280] = 0;
disk_mem[ 1281] = 0;
disk_mem[ 1282] = 0;
disk_mem[ 1283] = 0;
disk_mem[ 1284] = 0;
disk_mem[ 1285] = 0;
disk_mem[ 1286] = 0;
disk_mem[ 1287] = 0;
disk_mem[ 1288] = 0;
disk_mem[ 1289] = 0;
disk_mem[ 1290] = 0;
disk_mem[ 1291] = 0;
disk_mem[ 1292] = 0;
disk_mem[ 1293] = 0;
disk_mem[ 1294] = 0;
disk_mem[ 1295] = 0;
disk_mem[ 1296] = 0;
disk_mem[ 1297] = 0;
disk_mem[ 1298] = 0;
disk_mem[ 1299] = 0;
disk_mem[ 1300] = 0;
disk_mem[ 1301] = 0;
disk_mem[ 1302] = 0;
disk_mem[ 1303] = 0;
disk_mem[ 1304] = 0;
disk_mem[ 1305] = 0;
disk_mem[ 1306] = 0;
disk_mem[ 1307] = 0;
disk_mem[ 1308] = 0;
disk_mem[ 1309] = 0;
disk_mem[ 1310] = 0;
disk_mem[ 1311] = 0;
disk_mem[ 1312] = 0;
disk_mem[ 1313] = 0;
disk_mem[ 1314] = 0;
disk_mem[ 1315] = 0;
disk_mem[ 1316] = 0;
disk_mem[ 1317] = 0;
disk_mem[ 1318] = 0;
disk_mem[ 1319] = 0;
disk_mem[ 1320] = 0;
disk_mem[ 1321] = 0;
disk_mem[ 1322] = 0;
disk_mem[ 1323] = 0;
disk_mem[ 1324] = 0;
disk_mem[ 1325] = 0;
disk_mem[ 1326] = 0;
disk_mem[ 1327] = 0;
disk_mem[ 1328] = 0;
disk_mem[ 1329] = 0;
disk_mem[ 1330] = 0;
disk_mem[ 1331] = 0;
disk_mem[ 1332] = 0;
disk_mem[ 1333] = 0;
disk_mem[ 1334] = 0;
disk_mem[ 1335] = 0;
disk_mem[ 1336] = 0;
disk_mem[ 1337] = 0;
disk_mem[ 1338] = 0;
disk_mem[ 1339] = 0;
disk_mem[ 1340] = 0;
disk_mem[ 1341] = 0;
disk_mem[ 1342] = 0;
disk_mem[ 1343] = 0;
disk_mem[ 1344] = 0;
disk_mem[ 1345] = 0;
disk_mem[ 1346] = 0;
disk_mem[ 1347] = 0;
disk_mem[ 1348] = 0;
disk_mem[ 1349] = 0;
disk_mem[ 1350] = 0;
disk_mem[ 1351] = 0;
disk_mem[ 1352] = 0;
disk_mem[ 1353] = 0;
disk_mem[ 1354] = 0;
disk_mem[ 1355] = 0;
disk_mem[ 1356] = 0;
disk_mem[ 1357] = 0;
disk_mem[ 1358] = 0;
disk_mem[ 1359] = 0;
disk_mem[ 1360] = 0;
disk_mem[ 1361] = 0;
disk_mem[ 1362] = 0;
disk_mem[ 1363] = 0;
disk_mem[ 1364] = 0;
disk_mem[ 1365] = 0;
disk_mem[ 1366] = 0;
disk_mem[ 1367] = 0;
disk_mem[ 1368] = 0;
disk_mem[ 1369] = 0;
disk_mem[ 1370] = 0;
disk_mem[ 1371] = 0;
disk_mem[ 1372] = 0;
disk_mem[ 1373] = 0;
disk_mem[ 1374] = 0;
disk_mem[ 1375] = 0;
disk_mem[ 1376] = 0;
disk_mem[ 1377] = 0;
disk_mem[ 1378] = 0;
disk_mem[ 1379] = 0;
disk_mem[ 1380] = 0;
disk_mem[ 1381] = 0;
disk_mem[ 1382] = 0;
disk_mem[ 1383] = 0;
disk_mem[ 1384] = 0;
disk_mem[ 1385] = 0;
disk_mem[ 1386] = 0;
disk_mem[ 1387] = 0;
disk_mem[ 1388] = 0;
disk_mem[ 1389] = 0;
disk_mem[ 1390] = 0;
disk_mem[ 1391] = 0;
disk_mem[ 1392] = 0;
disk_mem[ 1393] = 0;
disk_mem[ 1394] = 0;
disk_mem[ 1395] = 0;
disk_mem[ 1396] = 0;
disk_mem[ 1397] = 0;
disk_mem[ 1398] = 0;
disk_mem[ 1399] = 0;
disk_mem[ 1400] = 0;
disk_mem[ 1401] = 0;
disk_mem[ 1402] = 0;
disk_mem[ 1403] = 0;
disk_mem[ 1404] = 0;
disk_mem[ 1405] = 0;
disk_mem[ 1406] = 0;
disk_mem[ 1407] = 0;
disk_mem[ 1408] = 0;
disk_mem[ 1409] = 0;
disk_mem[ 1410] = 0;
disk_mem[ 1411] = 0;
disk_mem[ 1412] = 0;
disk_mem[ 1413] = 0;
disk_mem[ 1414] = 0;
disk_mem[ 1415] = 0;
disk_mem[ 1416] = 0;
disk_mem[ 1417] = 0;
disk_mem[ 1418] = 0;
disk_mem[ 1419] = 0;
disk_mem[ 1420] = 0;
disk_mem[ 1421] = 0;
disk_mem[ 1422] = 0;
disk_mem[ 1423] = 0;
disk_mem[ 1424] = 0;
disk_mem[ 1425] = 0;
disk_mem[ 1426] = 0;
disk_mem[ 1427] = 0;
disk_mem[ 1428] = 0;
disk_mem[ 1429] = 0;
disk_mem[ 1430] = 0;
disk_mem[ 1431] = 0;
disk_mem[ 1432] = 0;
disk_mem[ 1433] = 0;
disk_mem[ 1434] = 0;
disk_mem[ 1435] = 0;
disk_mem[ 1436] = 0;
disk_mem[ 1437] = 0;
disk_mem[ 1438] = 0;
disk_mem[ 1439] = 0;
disk_mem[ 1440] = 0;
disk_mem[ 1441] = 0;
disk_mem[ 1442] = 0;
disk_mem[ 1443] = 0;
disk_mem[ 1444] = 0;
disk_mem[ 1445] = 0;
disk_mem[ 1446] = 0;
disk_mem[ 1447] = 0;
disk_mem[ 1448] = 0;
disk_mem[ 1449] = 0;
disk_mem[ 1450] = 0;
disk_mem[ 1451] = 0;
disk_mem[ 1452] = 0;
disk_mem[ 1453] = 0;
disk_mem[ 1454] = 0;
disk_mem[ 1455] = 0;
disk_mem[ 1456] = 0;
disk_mem[ 1457] = 0;
disk_mem[ 1458] = 0;
disk_mem[ 1459] = 0;
disk_mem[ 1460] = 0;
disk_mem[ 1461] = 0;
disk_mem[ 1462] = 0;
disk_mem[ 1463] = 0;
disk_mem[ 1464] = 0;
disk_mem[ 1465] = 0;
disk_mem[ 1466] = 0;
disk_mem[ 1467] = 0;
disk_mem[ 1468] = 0;
disk_mem[ 1469] = 0;
disk_mem[ 1470] = 0;
disk_mem[ 1471] = 0;
disk_mem[ 1472] = 0;
disk_mem[ 1473] = 0;
disk_mem[ 1474] = 0;
disk_mem[ 1475] = 0;
disk_mem[ 1476] = 0;
disk_mem[ 1477] = 0;
disk_mem[ 1478] = 0;
disk_mem[ 1479] = 0;
disk_mem[ 1480] = 0;
disk_mem[ 1481] = 0;
disk_mem[ 1482] = 0;
disk_mem[ 1483] = 0;
disk_mem[ 1484] = 0;
disk_mem[ 1485] = 0;
disk_mem[ 1486] = 0;
disk_mem[ 1487] = 0;
disk_mem[ 1488] = 0;
disk_mem[ 1489] = 0;
disk_mem[ 1490] = 0;
disk_mem[ 1491] = 0;
disk_mem[ 1492] = 0;
disk_mem[ 1493] = 0;
disk_mem[ 1494] = 0;
disk_mem[ 1495] = 0;
disk_mem[ 1496] = 0;
disk_mem[ 1497] = 0;
disk_mem[ 1498] = 0;
disk_mem[ 1499] = 0;
disk_mem[ 1500] = 0;
disk_mem[ 1501] = 0;
disk_mem[ 1502] = 0;
disk_mem[ 1503] = 0;
disk_mem[ 1504] = 0;
disk_mem[ 1505] = 0;
disk_mem[ 1506] = 0;
disk_mem[ 1507] = 0;
disk_mem[ 1508] = 0;
disk_mem[ 1509] = 0;
disk_mem[ 1510] = 0;
disk_mem[ 1511] = 0;
disk_mem[ 1512] = 0;
disk_mem[ 1513] = 0;
disk_mem[ 1514] = 0;
disk_mem[ 1515] = 0;
disk_mem[ 1516] = 0;
disk_mem[ 1517] = 0;
disk_mem[ 1518] = 0;
disk_mem[ 1519] = 0;
disk_mem[ 1520] = 0;
disk_mem[ 1521] = 0;
disk_mem[ 1522] = 0;
disk_mem[ 1523] = 0;
disk_mem[ 1524] = 0;
disk_mem[ 1525] = 0;
disk_mem[ 1526] = 0;
disk_mem[ 1527] = 0;
disk_mem[ 1528] = 0;
disk_mem[ 1529] = 0;
disk_mem[ 1530] = 0;
disk_mem[ 1531] = 0;
disk_mem[ 1532] = 0;
disk_mem[ 1533] = 0;
disk_mem[ 1534] = 0;
disk_mem[ 1535] = 0;
disk_mem[ 1536] = 0;
disk_mem[ 1537] = 0;
disk_mem[ 1538] = 0;
disk_mem[ 1539] = 0;
disk_mem[ 1540] = 0;
disk_mem[ 1541] = 0;
disk_mem[ 1542] = 0;
disk_mem[ 1543] = 0;
disk_mem[ 1544] = 0;
disk_mem[ 1545] = 0;
disk_mem[ 1546] = 0;
disk_mem[ 1547] = 0;
disk_mem[ 1548] = 0;
disk_mem[ 1549] = 0;
disk_mem[ 1550] = 0;
disk_mem[ 1551] = 0;
disk_mem[ 1552] = 0;
disk_mem[ 1553] = 0;
disk_mem[ 1554] = 0;
disk_mem[ 1555] = 0;
disk_mem[ 1556] = 0;
disk_mem[ 1557] = 0;
disk_mem[ 1558] = 0;
disk_mem[ 1559] = 0;
disk_mem[ 1560] = 0;
disk_mem[ 1561] = 0;
disk_mem[ 1562] = 0;
disk_mem[ 1563] = 0;
disk_mem[ 1564] = 0;
disk_mem[ 1565] = 0;
disk_mem[ 1566] = 0;
disk_mem[ 1567] = 0;
disk_mem[ 1568] = 0;
disk_mem[ 1569] = 0;
disk_mem[ 1570] = 0;
disk_mem[ 1571] = 0;
disk_mem[ 1572] = 0;
disk_mem[ 1573] = 0;
disk_mem[ 1574] = 0;
disk_mem[ 1575] = 0;
disk_mem[ 1576] = 0;
disk_mem[ 1577] = 0;
disk_mem[ 1578] = 0;
disk_mem[ 1579] = 0;
disk_mem[ 1580] = 0;
disk_mem[ 1581] = 0;
disk_mem[ 1582] = 0;
disk_mem[ 1583] = 0;
disk_mem[ 1584] = 0;
disk_mem[ 1585] = 0;
disk_mem[ 1586] = 0;
disk_mem[ 1587] = 0;
disk_mem[ 1588] = 0;
disk_mem[ 1589] = 0;
disk_mem[ 1590] = 0;
disk_mem[ 1591] = 0;
disk_mem[ 1592] = 0;
disk_mem[ 1593] = 0;
disk_mem[ 1594] = 0;
disk_mem[ 1595] = 0;
disk_mem[ 1596] = 0;
disk_mem[ 1597] = 0;
disk_mem[ 1598] = 0;
disk_mem[ 1599] = 0;
disk_mem[ 1600] = 0;
disk_mem[ 1601] = 0;
disk_mem[ 1602] = 0;
disk_mem[ 1603] = 0;
disk_mem[ 1604] = 0;
disk_mem[ 1605] = 0;
disk_mem[ 1606] = 0;
disk_mem[ 1607] = 0;
disk_mem[ 1608] = 0;
disk_mem[ 1609] = 0;
disk_mem[ 1610] = 0;
disk_mem[ 1611] = 0;
disk_mem[ 1612] = 0;
disk_mem[ 1613] = 0;
disk_mem[ 1614] = 0;
disk_mem[ 1615] = 0;
disk_mem[ 1616] = 0;
disk_mem[ 1617] = 0;
disk_mem[ 1618] = 0;
disk_mem[ 1619] = 0;
disk_mem[ 1620] = 0;
disk_mem[ 1621] = 0;
disk_mem[ 1622] = 0;
disk_mem[ 1623] = 0;
disk_mem[ 1624] = 0;
disk_mem[ 1625] = 0;
disk_mem[ 1626] = 0;
disk_mem[ 1627] = 0;
disk_mem[ 1628] = 0;
disk_mem[ 1629] = 0;
disk_mem[ 1630] = 0;
disk_mem[ 1631] = 0;
disk_mem[ 1632] = 0;
disk_mem[ 1633] = 0;
disk_mem[ 1634] = 0;
disk_mem[ 1635] = 0;
disk_mem[ 1636] = 0;
disk_mem[ 1637] = 0;
disk_mem[ 1638] = 0;
disk_mem[ 1639] = 0;
disk_mem[ 1640] = 0;
disk_mem[ 1641] = 0;
disk_mem[ 1642] = 0;
disk_mem[ 1643] = 0;
disk_mem[ 1644] = 0;
disk_mem[ 1645] = 0;
disk_mem[ 1646] = 0;
disk_mem[ 1647] = 0;
disk_mem[ 1648] = 0;
disk_mem[ 1649] = 0;
disk_mem[ 1650] = 0;
disk_mem[ 1651] = 0;
disk_mem[ 1652] = 0;
disk_mem[ 1653] = 0;
disk_mem[ 1654] = 0;
disk_mem[ 1655] = 0;
disk_mem[ 1656] = 0;
disk_mem[ 1657] = 0;
disk_mem[ 1658] = 0;
disk_mem[ 1659] = 0;
disk_mem[ 1660] = 0;
disk_mem[ 1661] = 0;
disk_mem[ 1662] = 0;
disk_mem[ 1663] = 0;
disk_mem[ 1664] = 0;
disk_mem[ 1665] = 0;
disk_mem[ 1666] = 0;
disk_mem[ 1667] = 0;
disk_mem[ 1668] = 0;
disk_mem[ 1669] = 0;
disk_mem[ 1670] = 0;
disk_mem[ 1671] = 0;
disk_mem[ 1672] = 0;
disk_mem[ 1673] = 0;
disk_mem[ 1674] = 0;
disk_mem[ 1675] = 0;
disk_mem[ 1676] = 0;
disk_mem[ 1677] = 0;
disk_mem[ 1678] = 0;
disk_mem[ 1679] = 0;
disk_mem[ 1680] = 0;
disk_mem[ 1681] = 0;
disk_mem[ 1682] = 0;
disk_mem[ 1683] = 0;
disk_mem[ 1684] = 0;
disk_mem[ 1685] = 0;
disk_mem[ 1686] = 0;
disk_mem[ 1687] = 0;
disk_mem[ 1688] = 0;
disk_mem[ 1689] = 0;
disk_mem[ 1690] = 0;
disk_mem[ 1691] = 0;
disk_mem[ 1692] = 0;
disk_mem[ 1693] = 0;
disk_mem[ 1694] = 0;
disk_mem[ 1695] = 0;
disk_mem[ 1696] = 0;
disk_mem[ 1697] = 0;
disk_mem[ 1698] = 0;
disk_mem[ 1699] = 0;
disk_mem[ 1700] = 0;
disk_mem[ 1701] = 0;
disk_mem[ 1702] = 0;
disk_mem[ 1703] = 0;
disk_mem[ 1704] = 0;
disk_mem[ 1705] = 0;
disk_mem[ 1706] = 0;
disk_mem[ 1707] = 0;
disk_mem[ 1708] = 0;
disk_mem[ 1709] = 0;
disk_mem[ 1710] = 0;
disk_mem[ 1711] = 0;
disk_mem[ 1712] = 0;
disk_mem[ 1713] = 0;
disk_mem[ 1714] = 0;
disk_mem[ 1715] = 0;
disk_mem[ 1716] = 0;
disk_mem[ 1717] = 0;
disk_mem[ 1718] = 0;
disk_mem[ 1719] = 0;
disk_mem[ 1720] = 0;
disk_mem[ 1721] = 0;
disk_mem[ 1722] = 0;
disk_mem[ 1723] = 0;
disk_mem[ 1724] = 0;
disk_mem[ 1725] = 0;
disk_mem[ 1726] = 0;
disk_mem[ 1727] = 0;
disk_mem[ 1728] = 0;
disk_mem[ 1729] = 0;
disk_mem[ 1730] = 0;
disk_mem[ 1731] = 0;
disk_mem[ 1732] = 0;
disk_mem[ 1733] = 0;
disk_mem[ 1734] = 0;
disk_mem[ 1735] = 0;
disk_mem[ 1736] = 0;
disk_mem[ 1737] = 0;
disk_mem[ 1738] = 0;
disk_mem[ 1739] = 0;
disk_mem[ 1740] = 0;
disk_mem[ 1741] = 0;
disk_mem[ 1742] = 0;
disk_mem[ 1743] = 0;
disk_mem[ 1744] = 0;
disk_mem[ 1745] = 0;
disk_mem[ 1746] = 0;
disk_mem[ 1747] = 0;
disk_mem[ 1748] = 0;
disk_mem[ 1749] = 0;
disk_mem[ 1750] = 0;
disk_mem[ 1751] = 0;
disk_mem[ 1752] = 0;
disk_mem[ 1753] = 0;
disk_mem[ 1754] = 0;
disk_mem[ 1755] = 0;
disk_mem[ 1756] = 0;
disk_mem[ 1757] = 0;
disk_mem[ 1758] = 0;
disk_mem[ 1759] = 0;
disk_mem[ 1760] = 0;
disk_mem[ 1761] = 0;
disk_mem[ 1762] = 0;
disk_mem[ 1763] = 0;
disk_mem[ 1764] = 0;
disk_mem[ 1765] = 0;
disk_mem[ 1766] = 0;
disk_mem[ 1767] = 0;
disk_mem[ 1768] = 0;
disk_mem[ 1769] = 0;
disk_mem[ 1770] = 0;
disk_mem[ 1771] = 0;
disk_mem[ 1772] = 0;
disk_mem[ 1773] = 0;
disk_mem[ 1774] = 0;
disk_mem[ 1775] = 0;
disk_mem[ 1776] = 0;
disk_mem[ 1777] = 0;
disk_mem[ 1778] = 0;
disk_mem[ 1779] = 0;
disk_mem[ 1780] = 0;
disk_mem[ 1781] = 0;
disk_mem[ 1782] = 0;
disk_mem[ 1783] = 0;
disk_mem[ 1784] = 0;
disk_mem[ 1785] = 0;
disk_mem[ 1786] = 0;
disk_mem[ 1787] = 0;
disk_mem[ 1788] = 0;
disk_mem[ 1789] = 0;
disk_mem[ 1790] = 0;
disk_mem[ 1791] = 0;
disk_mem[ 1792] = 0;
disk_mem[ 1793] = 0;
disk_mem[ 1794] = 0;
disk_mem[ 1795] = 0;
disk_mem[ 1796] = 0;
disk_mem[ 1797] = 0;
disk_mem[ 1798] = 0;
disk_mem[ 1799] = 0;
disk_mem[ 1800] = 0;
disk_mem[ 1801] = 0;
disk_mem[ 1802] = 0;
disk_mem[ 1803] = 0;
disk_mem[ 1804] = 0;
disk_mem[ 1805] = 0;
disk_mem[ 1806] = 0;
disk_mem[ 1807] = 0;
disk_mem[ 1808] = 0;
disk_mem[ 1809] = 0;
disk_mem[ 1810] = 0;
disk_mem[ 1811] = 0;
disk_mem[ 1812] = 0;
disk_mem[ 1813] = 0;
disk_mem[ 1814] = 0;
disk_mem[ 1815] = 0;
disk_mem[ 1816] = 0;
disk_mem[ 1817] = 0;
disk_mem[ 1818] = 0;
disk_mem[ 1819] = 0;
disk_mem[ 1820] = 0;
disk_mem[ 1821] = 0;
disk_mem[ 1822] = 0;
disk_mem[ 1823] = 0;
disk_mem[ 1824] = 0;
disk_mem[ 1825] = 0;
disk_mem[ 1826] = 0;
disk_mem[ 1827] = 0;
disk_mem[ 1828] = 0;
disk_mem[ 1829] = 0;
disk_mem[ 1830] = 0;
disk_mem[ 1831] = 0;
disk_mem[ 1832] = 0;
disk_mem[ 1833] = 0;
disk_mem[ 1834] = 0;
disk_mem[ 1835] = 0;
disk_mem[ 1836] = 0;
disk_mem[ 1837] = 0;
disk_mem[ 1838] = 0;
disk_mem[ 1839] = 0;
disk_mem[ 1840] = 0;
disk_mem[ 1841] = 0;
disk_mem[ 1842] = 0;
disk_mem[ 1843] = 0;
disk_mem[ 1844] = 0;
disk_mem[ 1845] = 0;
disk_mem[ 1846] = 0;
disk_mem[ 1847] = 0;
disk_mem[ 1848] = 0;
disk_mem[ 1849] = 0;
disk_mem[ 1850] = 0;
disk_mem[ 1851] = 0;
disk_mem[ 1852] = 0;
disk_mem[ 1853] = 0;
disk_mem[ 1854] = 0;
disk_mem[ 1855] = 0;
disk_mem[ 1856] = 0;
disk_mem[ 1857] = 0;
disk_mem[ 1858] = 0;
disk_mem[ 1859] = 0;
disk_mem[ 1860] = 0;
disk_mem[ 1861] = 0;
disk_mem[ 1862] = 0;
disk_mem[ 1863] = 0;
disk_mem[ 1864] = 0;
disk_mem[ 1865] = 0;
disk_mem[ 1866] = 0;
disk_mem[ 1867] = 0;
disk_mem[ 1868] = 0;
disk_mem[ 1869] = 0;
disk_mem[ 1870] = 0;
disk_mem[ 1871] = 0;
disk_mem[ 1872] = 0;
disk_mem[ 1873] = 0;
disk_mem[ 1874] = 0;
disk_mem[ 1875] = 0;
disk_mem[ 1876] = 0;
disk_mem[ 1877] = 0;
disk_mem[ 1878] = 0;
disk_mem[ 1879] = 0;
disk_mem[ 1880] = 0;
disk_mem[ 1881] = 0;
disk_mem[ 1882] = 0;
disk_mem[ 1883] = 0;
disk_mem[ 1884] = 0;
disk_mem[ 1885] = 0;
disk_mem[ 1886] = 0;
disk_mem[ 1887] = 0;
disk_mem[ 1888] = 0;
disk_mem[ 1889] = 0;
disk_mem[ 1890] = 0;
disk_mem[ 1891] = 0;
disk_mem[ 1892] = 0;
disk_mem[ 1893] = 0;
disk_mem[ 1894] = 0;
disk_mem[ 1895] = 0;
disk_mem[ 1896] = 0;
disk_mem[ 1897] = 0;
disk_mem[ 1898] = 0;
disk_mem[ 1899] = 0;
disk_mem[ 1900] = 0;
disk_mem[ 1901] = 0;
disk_mem[ 1902] = 0;
disk_mem[ 1903] = 0;
disk_mem[ 1904] = 0;
disk_mem[ 1905] = 0;
disk_mem[ 1906] = 0;
disk_mem[ 1907] = 0;
disk_mem[ 1908] = 0;
disk_mem[ 1909] = 0;
disk_mem[ 1910] = 0;
disk_mem[ 1911] = 0;
disk_mem[ 1912] = 0;
disk_mem[ 1913] = 0;
disk_mem[ 1914] = 0;
disk_mem[ 1915] = 0;
disk_mem[ 1916] = 0;
disk_mem[ 1917] = 0;
disk_mem[ 1918] = 0;
disk_mem[ 1919] = 0;
disk_mem[ 1920] = 0;
disk_mem[ 1921] = 0;
disk_mem[ 1922] = 0;
disk_mem[ 1923] = 0;
disk_mem[ 1924] = 0;
disk_mem[ 1925] = 0;
disk_mem[ 1926] = 0;
disk_mem[ 1927] = 0;
disk_mem[ 1928] = 0;
disk_mem[ 1929] = 0;
disk_mem[ 1930] = 0;
disk_mem[ 1931] = 0;
disk_mem[ 1932] = 0;
disk_mem[ 1933] = 0;
disk_mem[ 1934] = 0;
disk_mem[ 1935] = 0;
disk_mem[ 1936] = 0;
disk_mem[ 1937] = 0;
disk_mem[ 1938] = 0;
disk_mem[ 1939] = 0;
disk_mem[ 1940] = 0;
disk_mem[ 1941] = 0;
disk_mem[ 1942] = 0;
disk_mem[ 1943] = 0;
disk_mem[ 1944] = 0;
disk_mem[ 1945] = 0;
disk_mem[ 1946] = 0;
disk_mem[ 1947] = 0;
disk_mem[ 1948] = 0;
disk_mem[ 1949] = 0;
disk_mem[ 1950] = 0;
disk_mem[ 1951] = 0;
disk_mem[ 1952] = 0;
disk_mem[ 1953] = 0;
disk_mem[ 1954] = 0;
disk_mem[ 1955] = 0;
disk_mem[ 1956] = 0;
disk_mem[ 1957] = 0;
disk_mem[ 1958] = 0;
disk_mem[ 1959] = 0;
disk_mem[ 1960] = 0;
disk_mem[ 1961] = 0;
disk_mem[ 1962] = 0;
disk_mem[ 1963] = 0;
disk_mem[ 1964] = 0;
disk_mem[ 1965] = 0;
disk_mem[ 1966] = 0;
disk_mem[ 1967] = 0;
disk_mem[ 1968] = 0;
disk_mem[ 1969] = 0;
disk_mem[ 1970] = 0;
disk_mem[ 1971] = 0;
disk_mem[ 1972] = 0;
disk_mem[ 1973] = 0;
disk_mem[ 1974] = 0;
disk_mem[ 1975] = 0;
disk_mem[ 1976] = 0;
disk_mem[ 1977] = 0;
disk_mem[ 1978] = 0;
disk_mem[ 1979] = 0;
disk_mem[ 1980] = 0;
disk_mem[ 1981] = 0;
disk_mem[ 1982] = 0;
disk_mem[ 1983] = 0;
disk_mem[ 1984] = 0;
disk_mem[ 1985] = 0;
disk_mem[ 1986] = 0;
disk_mem[ 1987] = 0;
disk_mem[ 1988] = 0;
disk_mem[ 1989] = 0;
disk_mem[ 1990] = 0;
disk_mem[ 1991] = 0;
disk_mem[ 1992] = 0;
disk_mem[ 1993] = 0;
disk_mem[ 1994] = 0;
disk_mem[ 1995] = 0;
disk_mem[ 1996] = 0;
disk_mem[ 1997] = 0;
disk_mem[ 1998] = 0;
disk_mem[ 1999] = 0;
disk_mem[ 2000] = 0;
disk_mem[ 2001] = 0;
disk_mem[ 2002] = 0;
disk_mem[ 2003] = 0;
disk_mem[ 2004] = 0;
disk_mem[ 2005] = 0;
disk_mem[ 2006] = 0;
disk_mem[ 2007] = 0;
disk_mem[ 2008] = 0;
disk_mem[ 2009] = 0;
disk_mem[ 2010] = 0;
disk_mem[ 2011] = 0;
disk_mem[ 2012] = 0;
disk_mem[ 2013] = 0;
disk_mem[ 2014] = 0;
disk_mem[ 2015] = 0;
disk_mem[ 2016] = 0;
disk_mem[ 2017] = 0;
disk_mem[ 2018] = 0;
disk_mem[ 2019] = 0;
disk_mem[ 2020] = 0;
disk_mem[ 2021] = 0;
disk_mem[ 2022] = 0;
disk_mem[ 2023] = 0;
disk_mem[ 2024] = 0;
disk_mem[ 2025] = 0;
disk_mem[ 2026] = 0;
disk_mem[ 2027] = 0;
disk_mem[ 2028] = 0;
disk_mem[ 2029] = 0;
disk_mem[ 2030] = 0;
disk_mem[ 2031] = 0;
disk_mem[ 2032] = 0;
disk_mem[ 2033] = 0;
disk_mem[ 2034] = 0;
disk_mem[ 2035] = 0;
disk_mem[ 2036] = 0;
disk_mem[ 2037] = 0;
disk_mem[ 2038] = 0;
disk_mem[ 2039] = 0;
disk_mem[ 2040] = 0;
disk_mem[ 2041] = 0;
disk_mem[ 2042] = 0;
disk_mem[ 2043] = 0;
disk_mem[ 2044] = 0;
disk_mem[ 2045] = 0;
disk_mem[ 2046] = 0;
disk_mem[ 2047] = 0;
disk_mem[ 2048] = 0;
disk_mem[ 2049] = 0;
disk_mem[ 2050] = 0;
disk_mem[ 2051] = 0;
disk_mem[ 2052] = 0;
disk_mem[ 2053] = 0;
disk_mem[ 2054] = 0;
disk_mem[ 2055] = 0;
disk_mem[ 2056] = 0;
disk_mem[ 2057] = 0;
disk_mem[ 2058] = 0;
disk_mem[ 2059] = 0;
disk_mem[ 2060] = 0;
disk_mem[ 2061] = 0;
disk_mem[ 2062] = 0;
disk_mem[ 2063] = 0;
disk_mem[ 2064] = 0;
disk_mem[ 2065] = 0;
disk_mem[ 2066] = 0;
disk_mem[ 2067] = 0;
disk_mem[ 2068] = 0;
disk_mem[ 2069] = 0;
disk_mem[ 2070] = 0;
disk_mem[ 2071] = 0;
disk_mem[ 2072] = 0;
disk_mem[ 2073] = 0;
disk_mem[ 2074] = 0;
disk_mem[ 2075] = 0;
disk_mem[ 2076] = 0;
disk_mem[ 2077] = 0;
disk_mem[ 2078] = 0;
disk_mem[ 2079] = 0;
disk_mem[ 2080] = 0;
disk_mem[ 2081] = 0;
disk_mem[ 2082] = 0;
disk_mem[ 2083] = 0;
disk_mem[ 2084] = 0;
disk_mem[ 2085] = 0;
disk_mem[ 2086] = 0;
disk_mem[ 2087] = 0;
disk_mem[ 2088] = 0;
disk_mem[ 2089] = 0;
disk_mem[ 2090] = 0;
disk_mem[ 2091] = 0;
disk_mem[ 2092] = 0;
disk_mem[ 2093] = 0;
disk_mem[ 2094] = 0;
disk_mem[ 2095] = 0;
disk_mem[ 2096] = 0;
disk_mem[ 2097] = 0;
disk_mem[ 2098] = 0;
disk_mem[ 2099] = 0;
disk_mem[ 2100] = 0;
disk_mem[ 2101] = 0;
disk_mem[ 2102] = 0;
disk_mem[ 2103] = 0;
disk_mem[ 2104] = 0;
disk_mem[ 2105] = 0;
disk_mem[ 2106] = 0;
disk_mem[ 2107] = 0;
disk_mem[ 2108] = 0;
disk_mem[ 2109] = 0;
disk_mem[ 2110] = 0;
disk_mem[ 2111] = 0;
disk_mem[ 2112] = 0;
disk_mem[ 2113] = 0;
disk_mem[ 2114] = 0;
disk_mem[ 2115] = 0;
disk_mem[ 2116] = 0;
disk_mem[ 2117] = 0;
disk_mem[ 2118] = 0;
disk_mem[ 2119] = 0;
disk_mem[ 2120] = 0;
disk_mem[ 2121] = 0;
disk_mem[ 2122] = 0;
disk_mem[ 2123] = 0;
disk_mem[ 2124] = 0;
disk_mem[ 2125] = 0;
disk_mem[ 2126] = 0;
disk_mem[ 2127] = 0;
disk_mem[ 2128] = 0;
disk_mem[ 2129] = 0;
disk_mem[ 2130] = 0;
disk_mem[ 2131] = 0;
disk_mem[ 2132] = 0;
disk_mem[ 2133] = 0;
disk_mem[ 2134] = 0;
disk_mem[ 2135] = 0;
disk_mem[ 2136] = 0;
disk_mem[ 2137] = 0;
disk_mem[ 2138] = 0;
disk_mem[ 2139] = 0;
disk_mem[ 2140] = 0;
disk_mem[ 2141] = 0;
disk_mem[ 2142] = 0;
disk_mem[ 2143] = 0;
disk_mem[ 2144] = 0;
disk_mem[ 2145] = 0;
disk_mem[ 2146] = 0;
disk_mem[ 2147] = 0;
disk_mem[ 2148] = 0;
disk_mem[ 2149] = 0;
disk_mem[ 2150] = 0;
disk_mem[ 2151] = 0;
disk_mem[ 2152] = 0;
disk_mem[ 2153] = 0;
disk_mem[ 2154] = 0;
disk_mem[ 2155] = 0;
disk_mem[ 2156] = 0;
disk_mem[ 2157] = 0;
disk_mem[ 2158] = 0;
disk_mem[ 2159] = 0;
disk_mem[ 2160] = 0;
disk_mem[ 2161] = 0;
disk_mem[ 2162] = 0;
disk_mem[ 2163] = 0;
disk_mem[ 2164] = 0;
disk_mem[ 2165] = 0;
disk_mem[ 2166] = 0;
disk_mem[ 2167] = 0;
disk_mem[ 2168] = 0;
disk_mem[ 2169] = 0;
disk_mem[ 2170] = 0;
disk_mem[ 2171] = 0;
disk_mem[ 2172] = 0;
disk_mem[ 2173] = 0;
disk_mem[ 2174] = 0;
disk_mem[ 2175] = 0;
disk_mem[ 2176] = 0;
disk_mem[ 2177] = 0;
disk_mem[ 2178] = 0;
disk_mem[ 2179] = 0;
disk_mem[ 2180] = 0;
disk_mem[ 2181] = 0;
disk_mem[ 2182] = 0;
disk_mem[ 2183] = 0;
disk_mem[ 2184] = 0;
disk_mem[ 2185] = 0;
disk_mem[ 2186] = 0;
disk_mem[ 2187] = 0;
disk_mem[ 2188] = 0;
disk_mem[ 2189] = 0;
disk_mem[ 2190] = 0;
disk_mem[ 2191] = 0;
disk_mem[ 2192] = 0;
disk_mem[ 2193] = 0;
disk_mem[ 2194] = 0;
disk_mem[ 2195] = 0;
disk_mem[ 2196] = 0;
disk_mem[ 2197] = 0;
disk_mem[ 2198] = 0;
disk_mem[ 2199] = 0;
disk_mem[ 2200] = 0;
disk_mem[ 2201] = 0;
disk_mem[ 2202] = 0;
disk_mem[ 2203] = 0;
disk_mem[ 2204] = 0;
disk_mem[ 2205] = 0;
disk_mem[ 2206] = 0;
disk_mem[ 2207] = 0;
disk_mem[ 2208] = 0;
disk_mem[ 2209] = 0;
disk_mem[ 2210] = 0;
disk_mem[ 2211] = 0;
disk_mem[ 2212] = 0;
disk_mem[ 2213] = 0;
disk_mem[ 2214] = 0;
disk_mem[ 2215] = 0;
disk_mem[ 2216] = 0;
disk_mem[ 2217] = 0;
disk_mem[ 2218] = 0;
disk_mem[ 2219] = 0;
disk_mem[ 2220] = 0;
disk_mem[ 2221] = 0;
disk_mem[ 2222] = 0;
disk_mem[ 2223] = 0;
disk_mem[ 2224] = 0;
disk_mem[ 2225] = 0;
disk_mem[ 2226] = 0;
disk_mem[ 2227] = 0;
disk_mem[ 2228] = 0;
disk_mem[ 2229] = 0;
disk_mem[ 2230] = 0;
disk_mem[ 2231] = 0;
disk_mem[ 2232] = 0;
disk_mem[ 2233] = 0;
disk_mem[ 2234] = 0;
disk_mem[ 2235] = 0;
disk_mem[ 2236] = 0;
disk_mem[ 2237] = 0;
disk_mem[ 2238] = 0;
disk_mem[ 2239] = 0;
disk_mem[ 2240] = 0;
disk_mem[ 2241] = 0;
disk_mem[ 2242] = 0;
disk_mem[ 2243] = 0;
disk_mem[ 2244] = 0;
disk_mem[ 2245] = 0;
disk_mem[ 2246] = 0;
disk_mem[ 2247] = 0;
disk_mem[ 2248] = 0;
disk_mem[ 2249] = 0;
disk_mem[ 2250] = 0;
disk_mem[ 2251] = 0;
disk_mem[ 2252] = 0;
disk_mem[ 2253] = 0;
disk_mem[ 2254] = 0;
disk_mem[ 2255] = 0;
disk_mem[ 2256] = 0;
disk_mem[ 2257] = 0;
disk_mem[ 2258] = 0;
disk_mem[ 2259] = 0;
disk_mem[ 2260] = 0;
disk_mem[ 2261] = 0;
disk_mem[ 2262] = 0;
disk_mem[ 2263] = 0;
disk_mem[ 2264] = 0;
disk_mem[ 2265] = 0;
disk_mem[ 2266] = 0;
disk_mem[ 2267] = 0;
disk_mem[ 2268] = 0;
disk_mem[ 2269] = 0;
disk_mem[ 2270] = 0;
disk_mem[ 2271] = 0;
disk_mem[ 2272] = 0;
disk_mem[ 2273] = 0;
disk_mem[ 2274] = 0;
disk_mem[ 2275] = 0;
disk_mem[ 2276] = 0;
disk_mem[ 2277] = 0;
disk_mem[ 2278] = 0;
disk_mem[ 2279] = 0;
disk_mem[ 2280] = 0;
disk_mem[ 2281] = 0;
disk_mem[ 2282] = 0;
disk_mem[ 2283] = 0;
disk_mem[ 2284] = 0;
disk_mem[ 2285] = 0;
disk_mem[ 2286] = 0;
disk_mem[ 2287] = 0;
disk_mem[ 2288] = 0;
disk_mem[ 2289] = 0;
disk_mem[ 2290] = 0;
disk_mem[ 2291] = 0;
disk_mem[ 2292] = 0;
disk_mem[ 2293] = 0;
disk_mem[ 2294] = 0;
disk_mem[ 2295] = 0;
disk_mem[ 2296] = 0;
disk_mem[ 2297] = 0;
disk_mem[ 2298] = 0;
disk_mem[ 2299] = 0;
disk_mem[ 2300] = 0;
disk_mem[ 2301] = 0;
disk_mem[ 2302] = 0;
disk_mem[ 2303] = 0;
disk_mem[ 2304] = 0;
disk_mem[ 2305] = 0;
disk_mem[ 2306] = 0;
disk_mem[ 2307] = 0;
disk_mem[ 2308] = 0;
disk_mem[ 2309] = 0;
disk_mem[ 2310] = 0;
disk_mem[ 2311] = 0;
disk_mem[ 2312] = 0;
disk_mem[ 2313] = 0;
disk_mem[ 2314] = 0;
disk_mem[ 2315] = 0;
disk_mem[ 2316] = 0;
disk_mem[ 2317] = 0;
disk_mem[ 2318] = 0;
disk_mem[ 2319] = 0;
disk_mem[ 2320] = 0;
disk_mem[ 2321] = 0;
disk_mem[ 2322] = 0;
disk_mem[ 2323] = 0;
disk_mem[ 2324] = 0;
disk_mem[ 2325] = 0;
disk_mem[ 2326] = 0;
disk_mem[ 2327] = 0;
disk_mem[ 2328] = 0;
disk_mem[ 2329] = 0;
disk_mem[ 2330] = 0;
disk_mem[ 2331] = 0;
disk_mem[ 2332] = 0;
disk_mem[ 2333] = 0;
disk_mem[ 2334] = 0;
disk_mem[ 2335] = 0;
disk_mem[ 2336] = 0;
disk_mem[ 2337] = 0;
disk_mem[ 2338] = 0;
disk_mem[ 2339] = 0;
disk_mem[ 2340] = 0;
disk_mem[ 2341] = 0;
disk_mem[ 2342] = 0;
disk_mem[ 2343] = 0;
disk_mem[ 2344] = 0;
disk_mem[ 2345] = 0;
disk_mem[ 2346] = 0;
disk_mem[ 2347] = 0;
disk_mem[ 2348] = 0;
disk_mem[ 2349] = 0;
disk_mem[ 2350] = 0;
disk_mem[ 2351] = 0;
disk_mem[ 2352] = 0;
disk_mem[ 2353] = 0;
disk_mem[ 2354] = 0;
disk_mem[ 2355] = 0;
disk_mem[ 2356] = 0;
disk_mem[ 2357] = 0;
disk_mem[ 2358] = 0;
disk_mem[ 2359] = 0;
disk_mem[ 2360] = 0;
disk_mem[ 2361] = 0;
disk_mem[ 2362] = 0;
disk_mem[ 2363] = 0;
disk_mem[ 2364] = 0;
disk_mem[ 2365] = 0;
disk_mem[ 2366] = 0;
disk_mem[ 2367] = 0;
disk_mem[ 2368] = 0;
disk_mem[ 2369] = 0;
disk_mem[ 2370] = 0;
disk_mem[ 2371] = 0;
disk_mem[ 2372] = 0;
disk_mem[ 2373] = 0;
disk_mem[ 2374] = 0;
disk_mem[ 2375] = 0;
disk_mem[ 2376] = 0;
disk_mem[ 2377] = 0;
disk_mem[ 2378] = 0;
disk_mem[ 2379] = 0;
disk_mem[ 2380] = 0;
disk_mem[ 2381] = 0;
disk_mem[ 2382] = 0;
disk_mem[ 2383] = 0;
disk_mem[ 2384] = 0;
disk_mem[ 2385] = 0;
disk_mem[ 2386] = 0;
disk_mem[ 2387] = 0;
disk_mem[ 2388] = 0;
disk_mem[ 2389] = 0;
disk_mem[ 2390] = 0;
disk_mem[ 2391] = 0;
disk_mem[ 2392] = 0;
disk_mem[ 2393] = 0;
disk_mem[ 2394] = 0;
disk_mem[ 2395] = 0;
disk_mem[ 2396] = 0;
disk_mem[ 2397] = 0;
disk_mem[ 2398] = 0;
disk_mem[ 2399] = 0;
disk_mem[ 2400] = 0;
disk_mem[ 2401] = 0;
disk_mem[ 2402] = 0;
disk_mem[ 2403] = 0;
disk_mem[ 2404] = 0;
disk_mem[ 2405] = 0;
disk_mem[ 2406] = 0;
disk_mem[ 2407] = 0;
disk_mem[ 2408] = 0;
disk_mem[ 2409] = 0;
disk_mem[ 2410] = 0;
disk_mem[ 2411] = 0;
disk_mem[ 2412] = 0;
disk_mem[ 2413] = 0;
disk_mem[ 2414] = 0;
disk_mem[ 2415] = 0;
disk_mem[ 2416] = 0;
disk_mem[ 2417] = 0;
disk_mem[ 2418] = 0;
disk_mem[ 2419] = 0;
disk_mem[ 2420] = 0;
disk_mem[ 2421] = 0;
disk_mem[ 2422] = 0;
disk_mem[ 2423] = 0;
disk_mem[ 2424] = 0;
disk_mem[ 2425] = 0;
disk_mem[ 2426] = 0;
disk_mem[ 2427] = 0;
disk_mem[ 2428] = 0;
disk_mem[ 2429] = 0;
disk_mem[ 2430] = 0;
disk_mem[ 2431] = 0;
disk_mem[ 2432] = 0;
disk_mem[ 2433] = 0;
disk_mem[ 2434] = 0;
disk_mem[ 2435] = 0;
disk_mem[ 2436] = 0;
disk_mem[ 2437] = 0;
disk_mem[ 2438] = 0;
disk_mem[ 2439] = 0;
disk_mem[ 2440] = 0;
disk_mem[ 2441] = 0;
disk_mem[ 2442] = 0;
disk_mem[ 2443] = 0;
disk_mem[ 2444] = 0;
disk_mem[ 2445] = 0;
disk_mem[ 2446] = 0;
disk_mem[ 2447] = 0;
disk_mem[ 2448] = 0;
disk_mem[ 2449] = 0;
disk_mem[ 2450] = 0;
disk_mem[ 2451] = 0;
disk_mem[ 2452] = 0;
disk_mem[ 2453] = 0;
disk_mem[ 2454] = 0;
disk_mem[ 2455] = 0;
disk_mem[ 2456] = 0;
disk_mem[ 2457] = 0;
disk_mem[ 2458] = 0;
disk_mem[ 2459] = 0;
disk_mem[ 2460] = 0;
disk_mem[ 2461] = 0;
disk_mem[ 2462] = 0;
disk_mem[ 2463] = 0;
disk_mem[ 2464] = 0;
disk_mem[ 2465] = 0;
disk_mem[ 2466] = 0;
disk_mem[ 2467] = 0;
disk_mem[ 2468] = 0;
disk_mem[ 2469] = 0;
disk_mem[ 2470] = 0;
disk_mem[ 2471] = 0;
disk_mem[ 2472] = 0;
disk_mem[ 2473] = 0;
disk_mem[ 2474] = 0;
disk_mem[ 2475] = 0;
disk_mem[ 2476] = 0;
disk_mem[ 2477] = 0;
disk_mem[ 2478] = 0;
disk_mem[ 2479] = 0;
disk_mem[ 2480] = 0;
disk_mem[ 2481] = 0;
disk_mem[ 2482] = 0;
disk_mem[ 2483] = 0;
disk_mem[ 2484] = 0;
disk_mem[ 2485] = 0;
disk_mem[ 2486] = 0;
disk_mem[ 2487] = 0;
disk_mem[ 2488] = 0;
disk_mem[ 2489] = 0;
disk_mem[ 2490] = 0;
disk_mem[ 2491] = 0;
disk_mem[ 2492] = 0;
disk_mem[ 2493] = 0;
disk_mem[ 2494] = 0;
disk_mem[ 2495] = 0;
disk_mem[ 2496] = 0;
disk_mem[ 2497] = 0;
disk_mem[ 2498] = 0;
disk_mem[ 2499] = 0;
disk_mem[ 2500] = 0;
disk_mem[ 2501] = 0;
disk_mem[ 2502] = 0;
disk_mem[ 2503] = 0;
disk_mem[ 2504] = 0;
disk_mem[ 2505] = 0;
disk_mem[ 2506] = 0;
disk_mem[ 2507] = 0;
disk_mem[ 2508] = 0;
disk_mem[ 2509] = 0;
disk_mem[ 2510] = 0;
disk_mem[ 2511] = 0;
disk_mem[ 2512] = 0;
disk_mem[ 2513] = 0;
disk_mem[ 2514] = 0;
disk_mem[ 2515] = 0;
disk_mem[ 2516] = 0;
disk_mem[ 2517] = 0;
disk_mem[ 2518] = 0;
disk_mem[ 2519] = 0;
disk_mem[ 2520] = 0;
disk_mem[ 2521] = 0;
disk_mem[ 2522] = 0;
disk_mem[ 2523] = 0;
disk_mem[ 2524] = 0;
disk_mem[ 2525] = 0;
disk_mem[ 2526] = 0;
disk_mem[ 2527] = 0;
disk_mem[ 2528] = 0;
disk_mem[ 2529] = 0;
disk_mem[ 2530] = 0;
disk_mem[ 2531] = 0;
disk_mem[ 2532] = 0;
disk_mem[ 2533] = 0;
disk_mem[ 2534] = 0;
disk_mem[ 2535] = 0;
disk_mem[ 2536] = 0;
disk_mem[ 2537] = 0;
disk_mem[ 2538] = 0;
disk_mem[ 2539] = 0;
disk_mem[ 2540] = 0;
disk_mem[ 2541] = 0;
disk_mem[ 2542] = 0;
disk_mem[ 2543] = 0;
disk_mem[ 2544] = 0;
disk_mem[ 2545] = 0;
disk_mem[ 2546] = 0;
disk_mem[ 2547] = 0;
disk_mem[ 2548] = 0;
disk_mem[ 2549] = 0;
disk_mem[ 2550] = 0;
disk_mem[ 2551] = 0;
disk_mem[ 2552] = 0;
disk_mem[ 2553] = 0;
disk_mem[ 2554] = 0;
disk_mem[ 2555] = 0;
disk_mem[ 2556] = 0;
disk_mem[ 2557] = 0;
disk_mem[ 2558] = 0;
disk_mem[ 2559] = 0;
disk_mem[ 2560] = 0;
disk_mem[ 2561] = 0;
disk_mem[ 2562] = 0;
disk_mem[ 2563] = 0;
disk_mem[ 2564] = 0;
disk_mem[ 2565] = 0;
disk_mem[ 2566] = 0;
disk_mem[ 2567] = 0;
disk_mem[ 2568] = 0;
disk_mem[ 2569] = 0;
disk_mem[ 2570] = 0;
disk_mem[ 2571] = 0;
disk_mem[ 2572] = 0;
disk_mem[ 2573] = 0;
disk_mem[ 2574] = 0;
disk_mem[ 2575] = 0;
disk_mem[ 2576] = 0;
disk_mem[ 2577] = 0;
disk_mem[ 2578] = 0;
disk_mem[ 2579] = 0;
disk_mem[ 2580] = 0;
disk_mem[ 2581] = 0;
disk_mem[ 2582] = 0;
disk_mem[ 2583] = 0;
disk_mem[ 2584] = 0;
disk_mem[ 2585] = 0;
disk_mem[ 2586] = 0;
disk_mem[ 2587] = 0;
disk_mem[ 2588] = 0;
disk_mem[ 2589] = 0;
disk_mem[ 2590] = 0;
disk_mem[ 2591] = 0;
disk_mem[ 2592] = 0;
disk_mem[ 2593] = 0;
disk_mem[ 2594] = 0;
disk_mem[ 2595] = 0;
disk_mem[ 2596] = 0;
disk_mem[ 2597] = 0;
disk_mem[ 2598] = 0;
disk_mem[ 2599] = 0;
disk_mem[ 2600] = 0;
disk_mem[ 2601] = 0;
disk_mem[ 2602] = 0;
disk_mem[ 2603] = 0;
disk_mem[ 2604] = 0;
disk_mem[ 2605] = 0;
disk_mem[ 2606] = 0;
disk_mem[ 2607] = 0;
disk_mem[ 2608] = 0;
disk_mem[ 2609] = 0;
disk_mem[ 2610] = 0;
disk_mem[ 2611] = 0;
disk_mem[ 2612] = 0;
disk_mem[ 2613] = 0;
disk_mem[ 2614] = 0;
disk_mem[ 2615] = 0;
disk_mem[ 2616] = 0;
disk_mem[ 2617] = 0;
disk_mem[ 2618] = 0;
disk_mem[ 2619] = 0;
disk_mem[ 2620] = 0;
disk_mem[ 2621] = 0;
disk_mem[ 2622] = 0;
disk_mem[ 2623] = 0;
disk_mem[ 2624] = 0;
disk_mem[ 2625] = 0;
disk_mem[ 2626] = 0;
disk_mem[ 2627] = 0;
disk_mem[ 2628] = 0;
disk_mem[ 2629] = 0;
disk_mem[ 2630] = 0;
disk_mem[ 2631] = 0;
disk_mem[ 2632] = 0;
disk_mem[ 2633] = 0;
disk_mem[ 2634] = 0;
disk_mem[ 2635] = 0;
disk_mem[ 2636] = 0;
disk_mem[ 2637] = 0;
disk_mem[ 2638] = 0;
disk_mem[ 2639] = 0;
disk_mem[ 2640] = 0;
disk_mem[ 2641] = 0;
disk_mem[ 2642] = 0;
disk_mem[ 2643] = 0;
disk_mem[ 2644] = 0;
disk_mem[ 2645] = 0;
disk_mem[ 2646] = 0;
disk_mem[ 2647] = 0;
disk_mem[ 2648] = 0;
disk_mem[ 2649] = 0;
disk_mem[ 2650] = 0;
disk_mem[ 2651] = 0;
disk_mem[ 2652] = 0;
disk_mem[ 2653] = 0;
disk_mem[ 2654] = 0;
disk_mem[ 2655] = 0;
disk_mem[ 2656] = 0;
disk_mem[ 2657] = 0;
disk_mem[ 2658] = 0;
disk_mem[ 2659] = 0;
disk_mem[ 2660] = 0;
disk_mem[ 2661] = 0;
disk_mem[ 2662] = 0;
disk_mem[ 2663] = 0;
disk_mem[ 2664] = 0;
disk_mem[ 2665] = 0;
disk_mem[ 2666] = 0;
disk_mem[ 2667] = 0;
disk_mem[ 2668] = 0;
disk_mem[ 2669] = 0;
disk_mem[ 2670] = 0;
disk_mem[ 2671] = 0;
disk_mem[ 2672] = 0;
disk_mem[ 2673] = 0;
disk_mem[ 2674] = 0;
disk_mem[ 2675] = 0;
disk_mem[ 2676] = 0;
disk_mem[ 2677] = 0;
disk_mem[ 2678] = 0;
disk_mem[ 2679] = 0;
disk_mem[ 2680] = 0;
disk_mem[ 2681] = 0;
disk_mem[ 2682] = 0;
disk_mem[ 2683] = 0;
disk_mem[ 2684] = 0;
disk_mem[ 2685] = 0;
disk_mem[ 2686] = 0;
disk_mem[ 2687] = 0;
disk_mem[ 2688] = 0;
disk_mem[ 2689] = 0;
disk_mem[ 2690] = 0;
disk_mem[ 2691] = 0;
disk_mem[ 2692] = 0;
disk_mem[ 2693] = 0;
disk_mem[ 2694] = 0;
disk_mem[ 2695] = 0;
disk_mem[ 2696] = 0;
disk_mem[ 2697] = 0;
disk_mem[ 2698] = 0;
disk_mem[ 2699] = 0;
disk_mem[ 2700] = 0;
disk_mem[ 2701] = 0;
disk_mem[ 2702] = 0;
disk_mem[ 2703] = 0;
disk_mem[ 2704] = 0;
disk_mem[ 2705] = 0;
disk_mem[ 2706] = 0;
disk_mem[ 2707] = 0;
disk_mem[ 2708] = 0;
disk_mem[ 2709] = 0;
disk_mem[ 2710] = 0;
disk_mem[ 2711] = 0;
disk_mem[ 2712] = 0;
disk_mem[ 2713] = 0;
disk_mem[ 2714] = 0;
disk_mem[ 2715] = 0;
disk_mem[ 2716] = 0;
disk_mem[ 2717] = 0;
disk_mem[ 2718] = 0;
disk_mem[ 2719] = 0;
disk_mem[ 2720] = 0;
disk_mem[ 2721] = 0;
disk_mem[ 2722] = 0;
disk_mem[ 2723] = 0;
disk_mem[ 2724] = 0;
disk_mem[ 2725] = 0;
disk_mem[ 2726] = 0;
disk_mem[ 2727] = 0;
disk_mem[ 2728] = 0;
disk_mem[ 2729] = 0;
disk_mem[ 2730] = 0;
disk_mem[ 2731] = 0;
disk_mem[ 2732] = 0;
disk_mem[ 2733] = 0;
disk_mem[ 2734] = 0;
disk_mem[ 2735] = 0;
disk_mem[ 2736] = 0;
disk_mem[ 2737] = 0;
disk_mem[ 2738] = 0;
disk_mem[ 2739] = 0;
disk_mem[ 2740] = 0;
disk_mem[ 2741] = 0;
disk_mem[ 2742] = 0;
disk_mem[ 2743] = 0;
disk_mem[ 2744] = 0;
disk_mem[ 2745] = 0;
disk_mem[ 2746] = 0;
disk_mem[ 2747] = 0;
disk_mem[ 2748] = 0;
disk_mem[ 2749] = 0;
disk_mem[ 2750] = 0;
disk_mem[ 2751] = 0;
disk_mem[ 2752] = 0;
disk_mem[ 2753] = 0;
disk_mem[ 2754] = 0;
disk_mem[ 2755] = 0;
disk_mem[ 2756] = 0;
disk_mem[ 2757] = 0;
disk_mem[ 2758] = 0;
disk_mem[ 2759] = 0;
disk_mem[ 2760] = 0;
disk_mem[ 2761] = 0;
disk_mem[ 2762] = 0;
disk_mem[ 2763] = 0;
disk_mem[ 2764] = 0;
disk_mem[ 2765] = 0;
disk_mem[ 2766] = 0;
disk_mem[ 2767] = 0;
disk_mem[ 2768] = 0;
disk_mem[ 2769] = 0;
disk_mem[ 2770] = 0;
disk_mem[ 2771] = 0;
disk_mem[ 2772] = 0;
disk_mem[ 2773] = 0;
disk_mem[ 2774] = 0;
disk_mem[ 2775] = 0;
disk_mem[ 2776] = 0;
disk_mem[ 2777] = 0;
disk_mem[ 2778] = 0;
disk_mem[ 2779] = 0;
disk_mem[ 2780] = 0;
disk_mem[ 2781] = 0;
disk_mem[ 2782] = 0;
disk_mem[ 2783] = 0;
disk_mem[ 2784] = 0;
disk_mem[ 2785] = 0;
disk_mem[ 2786] = 0;
disk_mem[ 2787] = 0;
disk_mem[ 2788] = 0;
disk_mem[ 2789] = 0;
disk_mem[ 2790] = 0;
disk_mem[ 2791] = 0;
disk_mem[ 2792] = 0;
disk_mem[ 2793] = 0;
disk_mem[ 2794] = 0;
disk_mem[ 2795] = 0;
disk_mem[ 2796] = 0;
disk_mem[ 2797] = 0;
disk_mem[ 2798] = 0;
disk_mem[ 2799] = 0;
disk_mem[ 2800] = 0;
disk_mem[ 2801] = 0;
disk_mem[ 2802] = 0;
disk_mem[ 2803] = 0;
disk_mem[ 2804] = 0;
disk_mem[ 2805] = 0;
disk_mem[ 2806] = 0;
disk_mem[ 2807] = 0;
disk_mem[ 2808] = 0;
disk_mem[ 2809] = 0;
disk_mem[ 2810] = 0;
disk_mem[ 2811] = 0;
disk_mem[ 2812] = 0;
disk_mem[ 2813] = 0;
disk_mem[ 2814] = 0;
disk_mem[ 2815] = 0;
disk_mem[ 2816] = 0;
disk_mem[ 2817] = 0;
disk_mem[ 2818] = 0;
disk_mem[ 2819] = 0;
disk_mem[ 2820] = 0;
disk_mem[ 2821] = 0;
disk_mem[ 2822] = 0;
disk_mem[ 2823] = 0;
disk_mem[ 2824] = 0;
disk_mem[ 2825] = 0;
disk_mem[ 2826] = 0;
disk_mem[ 2827] = 0;
disk_mem[ 2828] = 0;
disk_mem[ 2829] = 0;
disk_mem[ 2830] = 0;
disk_mem[ 2831] = 0;
disk_mem[ 2832] = 0;
disk_mem[ 2833] = 0;
disk_mem[ 2834] = 0;
disk_mem[ 2835] = 0;
disk_mem[ 2836] = 0;
disk_mem[ 2837] = 0;
disk_mem[ 2838] = 0;
disk_mem[ 2839] = 0;
disk_mem[ 2840] = 0;
disk_mem[ 2841] = 0;
disk_mem[ 2842] = 0;
disk_mem[ 2843] = 0;
disk_mem[ 2844] = 0;
disk_mem[ 2845] = 0;
disk_mem[ 2846] = 0;
disk_mem[ 2847] = 0;
disk_mem[ 2848] = 0;
disk_mem[ 2849] = 0;
disk_mem[ 2850] = 0;
disk_mem[ 2851] = 0;
disk_mem[ 2852] = 0;
disk_mem[ 2853] = 0;
disk_mem[ 2854] = 0;
disk_mem[ 2855] = 0;
disk_mem[ 2856] = 0;
disk_mem[ 2857] = 0;
disk_mem[ 2858] = 0;
disk_mem[ 2859] = 0;
disk_mem[ 2860] = 0;
disk_mem[ 2861] = 0;
disk_mem[ 2862] = 0;
disk_mem[ 2863] = 0;
disk_mem[ 2864] = 0;
disk_mem[ 2865] = 0;
disk_mem[ 2866] = 0;
disk_mem[ 2867] = 0;
disk_mem[ 2868] = 0;
disk_mem[ 2869] = 0;
disk_mem[ 2870] = 0;
disk_mem[ 2871] = 0;
disk_mem[ 2872] = 0;
disk_mem[ 2873] = 0;
disk_mem[ 2874] = 0;
disk_mem[ 2875] = 0;
disk_mem[ 2876] = 0;
disk_mem[ 2877] = 0;
disk_mem[ 2878] = 0;
disk_mem[ 2879] = 0;
disk_mem[ 2880] = 0;
disk_mem[ 2881] = 0;
disk_mem[ 2882] = 0;
disk_mem[ 2883] = 0;
disk_mem[ 2884] = 0;
disk_mem[ 2885] = 0;
disk_mem[ 2886] = 0;
disk_mem[ 2887] = 0;
disk_mem[ 2888] = 0;
disk_mem[ 2889] = 0;
disk_mem[ 2890] = 0;
disk_mem[ 2891] = 0;
disk_mem[ 2892] = 0;
disk_mem[ 2893] = 0;
disk_mem[ 2894] = 0;
disk_mem[ 2895] = 0;
disk_mem[ 2896] = 0;
disk_mem[ 2897] = 0;
disk_mem[ 2898] = 0;
disk_mem[ 2899] = 0;
disk_mem[ 2900] = 0;
disk_mem[ 2901] = 0;
disk_mem[ 2902] = 0;
disk_mem[ 2903] = 0;
disk_mem[ 2904] = 0;
disk_mem[ 2905] = 0;
disk_mem[ 2906] = 0;
disk_mem[ 2907] = 0;
disk_mem[ 2908] = 0;
disk_mem[ 2909] = 0;
disk_mem[ 2910] = 0;
disk_mem[ 2911] = 0;
disk_mem[ 2912] = 0;
disk_mem[ 2913] = 0;
disk_mem[ 2914] = 0;
disk_mem[ 2915] = 0;
disk_mem[ 2916] = 0;
disk_mem[ 2917] = 0;
disk_mem[ 2918] = 0;
disk_mem[ 2919] = 0;
disk_mem[ 2920] = 0;
disk_mem[ 2921] = 0;
disk_mem[ 2922] = 0;
disk_mem[ 2923] = 0;
disk_mem[ 2924] = 0;
disk_mem[ 2925] = 0;
disk_mem[ 2926] = 0;
disk_mem[ 2927] = 0;
disk_mem[ 2928] = 0;
disk_mem[ 2929] = 0;
disk_mem[ 2930] = 0;
disk_mem[ 2931] = 0;
disk_mem[ 2932] = 0;
disk_mem[ 2933] = 0;
disk_mem[ 2934] = 0;
disk_mem[ 2935] = 0;
disk_mem[ 2936] = 0;
disk_mem[ 2937] = 0;
disk_mem[ 2938] = 0;
disk_mem[ 2939] = 0;
disk_mem[ 2940] = 0;
disk_mem[ 2941] = 0;
disk_mem[ 2942] = 0;
disk_mem[ 2943] = 0;
disk_mem[ 2944] = 0;
disk_mem[ 2945] = 0;
disk_mem[ 2946] = 0;
disk_mem[ 2947] = 0;
disk_mem[ 2948] = 0;
disk_mem[ 2949] = 0;
disk_mem[ 2950] = 0;
disk_mem[ 2951] = 0;
disk_mem[ 2952] = 0;
disk_mem[ 2953] = 0;
disk_mem[ 2954] = 0;
disk_mem[ 2955] = 0;
disk_mem[ 2956] = 0;
disk_mem[ 2957] = 0;
disk_mem[ 2958] = 0;
disk_mem[ 2959] = 0;
disk_mem[ 2960] = 0;
disk_mem[ 2961] = 0;
disk_mem[ 2962] = 0;
disk_mem[ 2963] = 0;
disk_mem[ 2964] = 0;
disk_mem[ 2965] = 0;
disk_mem[ 2966] = 0;
disk_mem[ 2967] = 0;
disk_mem[ 2968] = 0;
disk_mem[ 2969] = 0;
disk_mem[ 2970] = 0;
disk_mem[ 2971] = 0;
disk_mem[ 2972] = 0;
disk_mem[ 2973] = 0;
disk_mem[ 2974] = 0;
disk_mem[ 2975] = 0;
disk_mem[ 2976] = 0;
disk_mem[ 2977] = 0;
disk_mem[ 2978] = 0;
disk_mem[ 2979] = 0;
disk_mem[ 2980] = 0;
disk_mem[ 2981] = 0;
disk_mem[ 2982] = 0;
disk_mem[ 2983] = 0;
disk_mem[ 2984] = 0;
disk_mem[ 2985] = 0;
disk_mem[ 2986] = 0;
disk_mem[ 2987] = 0;
disk_mem[ 2988] = 0;
disk_mem[ 2989] = 0;
disk_mem[ 2990] = 0;
disk_mem[ 2991] = 0;
disk_mem[ 2992] = 0;
disk_mem[ 2993] = 0;
disk_mem[ 2994] = 0;
disk_mem[ 2995] = 0;
disk_mem[ 2996] = 0;
disk_mem[ 2997] = 0;
disk_mem[ 2998] = 0;
disk_mem[ 2999] = 0;
disk_mem[ 3000] = 0;
disk_mem[ 3001] = 0;
disk_mem[ 3002] = 0;
disk_mem[ 3003] = 0;
disk_mem[ 3004] = 0;
disk_mem[ 3005] = 0;
disk_mem[ 3006] = 0;
disk_mem[ 3007] = 0;
disk_mem[ 3008] = 0;
disk_mem[ 3009] = 0;
disk_mem[ 3010] = 0;
disk_mem[ 3011] = 0;
disk_mem[ 3012] = 0;
disk_mem[ 3013] = 0;
disk_mem[ 3014] = 0;
disk_mem[ 3015] = 0;
disk_mem[ 3016] = 0;
disk_mem[ 3017] = 0;
disk_mem[ 3018] = 0;
disk_mem[ 3019] = 0;
disk_mem[ 3020] = 0;
disk_mem[ 3021] = 0;
disk_mem[ 3022] = 0;
disk_mem[ 3023] = 0;
disk_mem[ 3024] = 0;
disk_mem[ 3025] = 0;
disk_mem[ 3026] = 0;
disk_mem[ 3027] = 0;
disk_mem[ 3028] = 0;
disk_mem[ 3029] = 0;
disk_mem[ 3030] = 0;
disk_mem[ 3031] = 0;
disk_mem[ 3032] = 0;
disk_mem[ 3033] = 0;
disk_mem[ 3034] = 0;
disk_mem[ 3035] = 0;
disk_mem[ 3036] = 0;
disk_mem[ 3037] = 0;
disk_mem[ 3038] = 0;
disk_mem[ 3039] = 0;
disk_mem[ 3040] = 0;
disk_mem[ 3041] = 0;
disk_mem[ 3042] = 0;
disk_mem[ 3043] = 0;
disk_mem[ 3044] = 0;
disk_mem[ 3045] = 0;
disk_mem[ 3046] = 0;
disk_mem[ 3047] = 0;
disk_mem[ 3048] = 0;
disk_mem[ 3049] = 0;
disk_mem[ 3050] = 0;
disk_mem[ 3051] = 0;
disk_mem[ 3052] = 0;
disk_mem[ 3053] = 0;
disk_mem[ 3054] = 0;
disk_mem[ 3055] = 0;
disk_mem[ 3056] = 0;
disk_mem[ 3057] = 0;
disk_mem[ 3058] = 0;
disk_mem[ 3059] = 0;
disk_mem[ 3060] = 0;
disk_mem[ 3061] = 0;
disk_mem[ 3062] = 0;
disk_mem[ 3063] = 0;
disk_mem[ 3064] = 0;
disk_mem[ 3065] = 0;
disk_mem[ 3066] = 0;
disk_mem[ 3067] = 0;
disk_mem[ 3068] = 0;
disk_mem[ 3069] = 0;
disk_mem[ 3070] = 0;
disk_mem[ 3071] = 0;
disk_mem[ 3072] = 0;
disk_mem[ 3073] = 0;
disk_mem[ 3074] = 0;
disk_mem[ 3075] = 0;
disk_mem[ 3076] = 0;
disk_mem[ 3077] = 0;
disk_mem[ 3078] = 0;
disk_mem[ 3079] = 0;
disk_mem[ 3080] = 0;
disk_mem[ 3081] = 0;
disk_mem[ 3082] = 0;
disk_mem[ 3083] = 0;
disk_mem[ 3084] = 0;
disk_mem[ 3085] = 0;
disk_mem[ 3086] = 0;
disk_mem[ 3087] = 0;
disk_mem[ 3088] = 0;
disk_mem[ 3089] = 0;
disk_mem[ 3090] = 0;
disk_mem[ 3091] = 0;
disk_mem[ 3092] = 0;
disk_mem[ 3093] = 0;
disk_mem[ 3094] = 0;
disk_mem[ 3095] = 0;
disk_mem[ 3096] = 0;
disk_mem[ 3097] = 0;
disk_mem[ 3098] = 0;
disk_mem[ 3099] = 0;
disk_mem[ 3100] = 0;
disk_mem[ 3101] = 0;
disk_mem[ 3102] = 0;
disk_mem[ 3103] = 0;
disk_mem[ 3104] = 0;
disk_mem[ 3105] = 0;
disk_mem[ 3106] = 0;
disk_mem[ 3107] = 0;
disk_mem[ 3108] = 0;
disk_mem[ 3109] = 0;
disk_mem[ 3110] = 0;
disk_mem[ 3111] = 0;
disk_mem[ 3112] = 0;
disk_mem[ 3113] = 0;
disk_mem[ 3114] = 0;
disk_mem[ 3115] = 0;
disk_mem[ 3116] = 0;
disk_mem[ 3117] = 0;
disk_mem[ 3118] = 0;
disk_mem[ 3119] = 0;
disk_mem[ 3120] = 0;
disk_mem[ 3121] = 0;
disk_mem[ 3122] = 0;
disk_mem[ 3123] = 0;
disk_mem[ 3124] = 0;
disk_mem[ 3125] = 0;
disk_mem[ 3126] = 0;
disk_mem[ 3127] = 0;
disk_mem[ 3128] = 0;
disk_mem[ 3129] = 0;
disk_mem[ 3130] = 0;
disk_mem[ 3131] = 0;
disk_mem[ 3132] = 0;
disk_mem[ 3133] = 0;
disk_mem[ 3134] = 0;
disk_mem[ 3135] = 0;
disk_mem[ 3136] = 0;
disk_mem[ 3137] = 0;
disk_mem[ 3138] = 0;
disk_mem[ 3139] = 0;
disk_mem[ 3140] = 0;
disk_mem[ 3141] = 0;
disk_mem[ 3142] = 0;
disk_mem[ 3143] = 0;
disk_mem[ 3144] = 0;
disk_mem[ 3145] = 0;
disk_mem[ 3146] = 0;
disk_mem[ 3147] = 0;
disk_mem[ 3148] = 0;
disk_mem[ 3149] = 0;
disk_mem[ 3150] = 0;
disk_mem[ 3151] = 0;
disk_mem[ 3152] = 0;
disk_mem[ 3153] = 0;
disk_mem[ 3154] = 0;
disk_mem[ 3155] = 0;
disk_mem[ 3156] = 0;
disk_mem[ 3157] = 0;
disk_mem[ 3158] = 0;
disk_mem[ 3159] = 0;
disk_mem[ 3160] = 0;
disk_mem[ 3161] = 0;
disk_mem[ 3162] = 0;
disk_mem[ 3163] = 0;
disk_mem[ 3164] = 0;
disk_mem[ 3165] = 0;
disk_mem[ 3166] = 0;
disk_mem[ 3167] = 0;
disk_mem[ 3168] = 0;
disk_mem[ 3169] = 0;
disk_mem[ 3170] = 0;
disk_mem[ 3171] = 0;
disk_mem[ 3172] = 0;
disk_mem[ 3173] = 0;
disk_mem[ 3174] = 0;
disk_mem[ 3175] = 0;
disk_mem[ 3176] = 0;
disk_mem[ 3177] = 0;
disk_mem[ 3178] = 0;
disk_mem[ 3179] = 0;
disk_mem[ 3180] = 0;
disk_mem[ 3181] = 0;
disk_mem[ 3182] = 0;
disk_mem[ 3183] = 0;
disk_mem[ 3184] = 0;
disk_mem[ 3185] = 0;
disk_mem[ 3186] = 0;
disk_mem[ 3187] = 0;
disk_mem[ 3188] = 0;
disk_mem[ 3189] = 0;
disk_mem[ 3190] = 0;
disk_mem[ 3191] = 0;
disk_mem[ 3192] = 0;
disk_mem[ 3193] = 0;
disk_mem[ 3194] = 0;
disk_mem[ 3195] = 0;
disk_mem[ 3196] = 0;
disk_mem[ 3197] = 0;
disk_mem[ 3198] = 0;
disk_mem[ 3199] = 0;
disk_mem[ 3200] = 0;
disk_mem[ 3201] = 0;
disk_mem[ 3202] = 0;
disk_mem[ 3203] = 0;
disk_mem[ 3204] = 0;
disk_mem[ 3205] = 0;
disk_mem[ 3206] = 0;
disk_mem[ 3207] = 0;
disk_mem[ 3208] = 0;
disk_mem[ 3209] = 0;
disk_mem[ 3210] = 0;
disk_mem[ 3211] = 0;
disk_mem[ 3212] = 0;
disk_mem[ 3213] = 0;
disk_mem[ 3214] = 0;
disk_mem[ 3215] = 0;
disk_mem[ 3216] = 0;
disk_mem[ 3217] = 0;
disk_mem[ 3218] = 0;
disk_mem[ 3219] = 0;
disk_mem[ 3220] = 0;
disk_mem[ 3221] = 0;
disk_mem[ 3222] = 0;
disk_mem[ 3223] = 0;
disk_mem[ 3224] = 0;
disk_mem[ 3225] = 0;
disk_mem[ 3226] = 0;
disk_mem[ 3227] = 0;
disk_mem[ 3228] = 0;
disk_mem[ 3229] = 0;
disk_mem[ 3230] = 0;
disk_mem[ 3231] = 0;
disk_mem[ 3232] = 0;
disk_mem[ 3233] = 0;
disk_mem[ 3234] = 0;
disk_mem[ 3235] = 0;
disk_mem[ 3236] = 0;
disk_mem[ 3237] = 0;
disk_mem[ 3238] = 0;
disk_mem[ 3239] = 0;
disk_mem[ 3240] = 0;
disk_mem[ 3241] = 0;
disk_mem[ 3242] = 0;
disk_mem[ 3243] = 0;
disk_mem[ 3244] = 0;
disk_mem[ 3245] = 0;
disk_mem[ 3246] = 0;
disk_mem[ 3247] = 0;
disk_mem[ 3248] = 0;
disk_mem[ 3249] = 0;
disk_mem[ 3250] = 0;
disk_mem[ 3251] = 0;
disk_mem[ 3252] = 0;
disk_mem[ 3253] = 0;
disk_mem[ 3254] = 0;
disk_mem[ 3255] = 0;
disk_mem[ 3256] = 0;
disk_mem[ 3257] = 0;
disk_mem[ 3258] = 0;
disk_mem[ 3259] = 0;
disk_mem[ 3260] = 0;
disk_mem[ 3261] = 0;
disk_mem[ 3262] = 0;
disk_mem[ 3263] = 0;
disk_mem[ 3264] = 0;
disk_mem[ 3265] = 0;
disk_mem[ 3266] = 0;
disk_mem[ 3267] = 0;
disk_mem[ 3268] = 0;
disk_mem[ 3269] = 0;
disk_mem[ 3270] = 0;
disk_mem[ 3271] = 0;
disk_mem[ 3272] = 0;
disk_mem[ 3273] = 0;
disk_mem[ 3274] = 0;
disk_mem[ 3275] = 0;
disk_mem[ 3276] = 0;
disk_mem[ 3277] = 0;
disk_mem[ 3278] = 0;
disk_mem[ 3279] = 0;
disk_mem[ 3280] = 0;
disk_mem[ 3281] = 0;
disk_mem[ 3282] = 0;
disk_mem[ 3283] = 0;
disk_mem[ 3284] = 0;
disk_mem[ 3285] = 0;
disk_mem[ 3286] = 0;
disk_mem[ 3287] = 0;
disk_mem[ 3288] = 0;
disk_mem[ 3289] = 0;
disk_mem[ 3290] = 0;
disk_mem[ 3291] = 0;
disk_mem[ 3292] = 0;
disk_mem[ 3293] = 0;
disk_mem[ 3294] = 0;
disk_mem[ 3295] = 0;
disk_mem[ 3296] = 0;
disk_mem[ 3297] = 0;
disk_mem[ 3298] = 0;
disk_mem[ 3299] = 0;
disk_mem[ 3300] = 0;
disk_mem[ 3301] = 0;
disk_mem[ 3302] = 0;
disk_mem[ 3303] = 0;
disk_mem[ 3304] = 0;
disk_mem[ 3305] = 0;
disk_mem[ 3306] = 0;
disk_mem[ 3307] = 0;
disk_mem[ 3308] = 0;
disk_mem[ 3309] = 0;
disk_mem[ 3310] = 0;
disk_mem[ 3311] = 0;
disk_mem[ 3312] = 0;
disk_mem[ 3313] = 0;
disk_mem[ 3314] = 0;
disk_mem[ 3315] = 0;
disk_mem[ 3316] = 0;
disk_mem[ 3317] = 0;
disk_mem[ 3318] = 0;
disk_mem[ 3319] = 0;
disk_mem[ 3320] = 0;
disk_mem[ 3321] = 0;
disk_mem[ 3322] = 0;
disk_mem[ 3323] = 0;
disk_mem[ 3324] = 0;
disk_mem[ 3325] = 0;
disk_mem[ 3326] = 0;
disk_mem[ 3327] = 0;
disk_mem[ 3328] = 0;
disk_mem[ 3329] = 0;
disk_mem[ 3330] = 0;
disk_mem[ 3331] = 0;
disk_mem[ 3332] = 0;
disk_mem[ 3333] = 0;
disk_mem[ 3334] = 0;
disk_mem[ 3335] = 0;
disk_mem[ 3336] = 0;
disk_mem[ 3337] = 0;
disk_mem[ 3338] = 0;
disk_mem[ 3339] = 0;
disk_mem[ 3340] = 0;
disk_mem[ 3341] = 0;
disk_mem[ 3342] = 0;
disk_mem[ 3343] = 0;
disk_mem[ 3344] = 0;
disk_mem[ 3345] = 0;
disk_mem[ 3346] = 0;
disk_mem[ 3347] = 0;
disk_mem[ 3348] = 0;
disk_mem[ 3349] = 0;
disk_mem[ 3350] = 0;
disk_mem[ 3351] = 0;
disk_mem[ 3352] = 0;
disk_mem[ 3353] = 0;
disk_mem[ 3354] = 0;
disk_mem[ 3355] = 0;
disk_mem[ 3356] = 0;
disk_mem[ 3357] = 0;
disk_mem[ 3358] = 0;
disk_mem[ 3359] = 0;
disk_mem[ 3360] = 0;
disk_mem[ 3361] = 0;
disk_mem[ 3362] = 0;
disk_mem[ 3363] = 0;
disk_mem[ 3364] = 0;
disk_mem[ 3365] = 0;
disk_mem[ 3366] = 0;
disk_mem[ 3367] = 0;
disk_mem[ 3368] = 0;
disk_mem[ 3369] = 0;
disk_mem[ 3370] = 0;
disk_mem[ 3371] = 0;
disk_mem[ 3372] = 0;
disk_mem[ 3373] = 0;
disk_mem[ 3374] = 0;
disk_mem[ 3375] = 0;
disk_mem[ 3376] = 0;
disk_mem[ 3377] = 0;
disk_mem[ 3378] = 0;
disk_mem[ 3379] = 0;
disk_mem[ 3380] = 0;
disk_mem[ 3381] = 0;
disk_mem[ 3382] = 0;
disk_mem[ 3383] = 0;
disk_mem[ 3384] = 0;
disk_mem[ 3385] = 0;
disk_mem[ 3386] = 0;
disk_mem[ 3387] = 0;
disk_mem[ 3388] = 0;
disk_mem[ 3389] = 0;
disk_mem[ 3390] = 0;
disk_mem[ 3391] = 0;
disk_mem[ 3392] = 0;
disk_mem[ 3393] = 0;
disk_mem[ 3394] = 0;
disk_mem[ 3395] = 0;
disk_mem[ 3396] = 0;
disk_mem[ 3397] = 0;
disk_mem[ 3398] = 0;
disk_mem[ 3399] = 0;
disk_mem[ 3400] = 0;
disk_mem[ 3401] = 0;
disk_mem[ 3402] = 0;
disk_mem[ 3403] = 0;
disk_mem[ 3404] = 0;
disk_mem[ 3405] = 0;
disk_mem[ 3406] = 0;
disk_mem[ 3407] = 0;
disk_mem[ 3408] = 0;
disk_mem[ 3409] = 0;
disk_mem[ 3410] = 0;
disk_mem[ 3411] = 0;
disk_mem[ 3412] = 0;
disk_mem[ 3413] = 0;
disk_mem[ 3414] = 0;
disk_mem[ 3415] = 0;
disk_mem[ 3416] = 0;
disk_mem[ 3417] = 0;
disk_mem[ 3418] = 0;
disk_mem[ 3419] = 0;
disk_mem[ 3420] = 0;
disk_mem[ 3421] = 0;
disk_mem[ 3422] = 0;
disk_mem[ 3423] = 0;
disk_mem[ 3424] = 0;
disk_mem[ 3425] = 0;
disk_mem[ 3426] = 0;
disk_mem[ 3427] = 0;
disk_mem[ 3428] = 0;
disk_mem[ 3429] = 0;
disk_mem[ 3430] = 0;
disk_mem[ 3431] = 0;
disk_mem[ 3432] = 0;
disk_mem[ 3433] = 0;
disk_mem[ 3434] = 0;
disk_mem[ 3435] = 0;
disk_mem[ 3436] = 0;
disk_mem[ 3437] = 0;
disk_mem[ 3438] = 0;
disk_mem[ 3439] = 0;
disk_mem[ 3440] = 0;
disk_mem[ 3441] = 0;
disk_mem[ 3442] = 0;
disk_mem[ 3443] = 0;
disk_mem[ 3444] = 0;
disk_mem[ 3445] = 0;
disk_mem[ 3446] = 0;
disk_mem[ 3447] = 0;
disk_mem[ 3448] = 0;
disk_mem[ 3449] = 0;
disk_mem[ 3450] = 0;
disk_mem[ 3451] = 0;
disk_mem[ 3452] = 0;
disk_mem[ 3453] = 0;
disk_mem[ 3454] = 0;
disk_mem[ 3455] = 0;
disk_mem[ 3456] = 0;
disk_mem[ 3457] = 0;
disk_mem[ 3458] = 0;
disk_mem[ 3459] = 0;
disk_mem[ 3460] = 0;
disk_mem[ 3461] = 0;
disk_mem[ 3462] = 0;
disk_mem[ 3463] = 0;
disk_mem[ 3464] = 0;
disk_mem[ 3465] = 0;
disk_mem[ 3466] = 0;
disk_mem[ 3467] = 0;
disk_mem[ 3468] = 0;
disk_mem[ 3469] = 0;
disk_mem[ 3470] = 0;
disk_mem[ 3471] = 0;
disk_mem[ 3472] = 0;
disk_mem[ 3473] = 0;
disk_mem[ 3474] = 0;
disk_mem[ 3475] = 0;
disk_mem[ 3476] = 0;
disk_mem[ 3477] = 0;
disk_mem[ 3478] = 0;
disk_mem[ 3479] = 0;
disk_mem[ 3480] = 0;
disk_mem[ 3481] = 0;
disk_mem[ 3482] = 0;
disk_mem[ 3483] = 0;
disk_mem[ 3484] = 0;
disk_mem[ 3485] = 0;
disk_mem[ 3486] = 0;
disk_mem[ 3487] = 0;
disk_mem[ 3488] = 0;
disk_mem[ 3489] = 0;
disk_mem[ 3490] = 0;
disk_mem[ 3491] = 0;
disk_mem[ 3492] = 0;
disk_mem[ 3493] = 0;
disk_mem[ 3494] = 0;
disk_mem[ 3495] = 0;
disk_mem[ 3496] = 0;
disk_mem[ 3497] = 0;
disk_mem[ 3498] = 0;
disk_mem[ 3499] = 0;
disk_mem[ 3500] = 0;
disk_mem[ 3501] = 0;
disk_mem[ 3502] = 0;
disk_mem[ 3503] = 0;
disk_mem[ 3504] = 0;
disk_mem[ 3505] = 0;
disk_mem[ 3506] = 0;
disk_mem[ 3507] = 0;
disk_mem[ 3508] = 0;
disk_mem[ 3509] = 0;
disk_mem[ 3510] = 0;
disk_mem[ 3511] = 0;
disk_mem[ 3512] = 0;
disk_mem[ 3513] = 0;
disk_mem[ 3514] = 0;
disk_mem[ 3515] = 0;
disk_mem[ 3516] = 0;
disk_mem[ 3517] = 0;
disk_mem[ 3518] = 0;
disk_mem[ 3519] = 0;
disk_mem[ 3520] = 0;
disk_mem[ 3521] = 0;
disk_mem[ 3522] = 0;
disk_mem[ 3523] = 0;
disk_mem[ 3524] = 0;
disk_mem[ 3525] = 0;
disk_mem[ 3526] = 0;
disk_mem[ 3527] = 0;
disk_mem[ 3528] = 0;
disk_mem[ 3529] = 0;
disk_mem[ 3530] = 0;
disk_mem[ 3531] = 0;
disk_mem[ 3532] = 0;
disk_mem[ 3533] = 0;
disk_mem[ 3534] = 0;
disk_mem[ 3535] = 0;
disk_mem[ 3536] = 0;
disk_mem[ 3537] = 0;
disk_mem[ 3538] = 0;
disk_mem[ 3539] = 0;
disk_mem[ 3540] = 0;
disk_mem[ 3541] = 0;
disk_mem[ 3542] = 0;
disk_mem[ 3543] = 0;
disk_mem[ 3544] = 0;
disk_mem[ 3545] = 0;
disk_mem[ 3546] = 0;
disk_mem[ 3547] = 0;
disk_mem[ 3548] = 0;
disk_mem[ 3549] = 0;
disk_mem[ 3550] = 0;
disk_mem[ 3551] = 0;
disk_mem[ 3552] = 0;
disk_mem[ 3553] = 0;
disk_mem[ 3554] = 0;
disk_mem[ 3555] = 0;
disk_mem[ 3556] = 0;
disk_mem[ 3557] = 0;
disk_mem[ 3558] = 0;
disk_mem[ 3559] = 0;
disk_mem[ 3560] = 0;
disk_mem[ 3561] = 0;
disk_mem[ 3562] = 0;
disk_mem[ 3563] = 0;
disk_mem[ 3564] = 0;
disk_mem[ 3565] = 0;
disk_mem[ 3566] = 0;
disk_mem[ 3567] = 0;
disk_mem[ 3568] = 0;
disk_mem[ 3569] = 0;
disk_mem[ 3570] = 0;
disk_mem[ 3571] = 0;
disk_mem[ 3572] = 0;
disk_mem[ 3573] = 0;
disk_mem[ 3574] = 0;
disk_mem[ 3575] = 0;
disk_mem[ 3576] = 0;
disk_mem[ 3577] = 0;
disk_mem[ 3578] = 0;
disk_mem[ 3579] = 0;
disk_mem[ 3580] = 0;
disk_mem[ 3581] = 0;
disk_mem[ 3582] = 0;
disk_mem[ 3583] = 0;
disk_mem[ 3584] = 'hF8;
disk_mem[ 3585] = 'hFF;
disk_mem[ 3586] = 'hFF;
disk_mem[ 3587] = 'hFF;
disk_mem[ 3588] = 'hFF;
disk_mem[ 3589] = 'hFF;
disk_mem[ 3590] = 'hFF;
disk_mem[ 3591] = 'hFF;
disk_mem[ 3592] = 'hFF;
disk_mem[ 3593] = 0;
disk_mem[ 3594] = 0;
disk_mem[ 3595] = 0;
disk_mem[ 3596] = 0;
disk_mem[ 3597] = 0;
disk_mem[ 3598] = 0;
disk_mem[ 3599] = 0;
disk_mem[ 3600] = 0;
disk_mem[ 3601] = 0;
disk_mem[ 3602] = 0;
disk_mem[ 3603] = 0;
disk_mem[ 3604] = 0;
disk_mem[ 3605] = 0;
disk_mem[ 3606] = 0;
disk_mem[ 3607] = 0;
disk_mem[ 3608] = 0;
disk_mem[ 3609] = 0;
disk_mem[ 3610] = 0;
disk_mem[ 3611] = 0;
disk_mem[ 3612] = 0;
disk_mem[ 3613] = 0;
disk_mem[ 3614] = 0;
disk_mem[ 3615] = 0;
disk_mem[ 3616] = 0;
disk_mem[ 3617] = 0;
disk_mem[ 3618] = 0;
disk_mem[ 3619] = 0;
disk_mem[ 3620] = 0;
disk_mem[ 3621] = 0;
disk_mem[ 3622] = 0;
disk_mem[ 3623] = 0;
disk_mem[ 3624] = 0;
disk_mem[ 3625] = 0;
disk_mem[ 3626] = 0;
disk_mem[ 3627] = 0;
disk_mem[ 3628] = 0;
disk_mem[ 3629] = 0;
disk_mem[ 3630] = 0;
disk_mem[ 3631] = 0;
disk_mem[ 3632] = 0;
disk_mem[ 3633] = 0;
disk_mem[ 3634] = 0;
disk_mem[ 3635] = 0;
disk_mem[ 3636] = 0;
disk_mem[ 3637] = 0;
disk_mem[ 3638] = 0;
disk_mem[ 3639] = 0;
disk_mem[ 3640] = 0;
disk_mem[ 3641] = 0;
disk_mem[ 3642] = 0;
disk_mem[ 3643] = 0;
disk_mem[ 3644] = 0;
disk_mem[ 3645] = 0;
disk_mem[ 3646] = 0;
disk_mem[ 3647] = 0;
disk_mem[ 3648] = 0;
disk_mem[ 3649] = 0;
disk_mem[ 3650] = 0;
disk_mem[ 3651] = 0;
disk_mem[ 3652] = 0;
disk_mem[ 3653] = 0;
disk_mem[ 3654] = 0;
disk_mem[ 3655] = 0;
disk_mem[ 3656] = 0;
disk_mem[ 3657] = 0;
disk_mem[ 3658] = 0;
disk_mem[ 3659] = 0;
disk_mem[ 3660] = 0;
disk_mem[ 3661] = 0;
disk_mem[ 3662] = 0;
disk_mem[ 3663] = 0;
disk_mem[ 3664] = 0;
disk_mem[ 3665] = 0;
disk_mem[ 3666] = 0;
disk_mem[ 3667] = 0;
disk_mem[ 3668] = 0;
disk_mem[ 3669] = 0;
disk_mem[ 3670] = 0;
disk_mem[ 3671] = 0;
disk_mem[ 3672] = 0;
disk_mem[ 3673] = 0;
disk_mem[ 3674] = 0;
disk_mem[ 3675] = 0;
disk_mem[ 3676] = 0;
disk_mem[ 3677] = 0;
disk_mem[ 3678] = 0;
disk_mem[ 3679] = 0;
disk_mem[ 3680] = 0;
disk_mem[ 3681] = 0;
disk_mem[ 3682] = 0;
disk_mem[ 3683] = 0;
disk_mem[ 3684] = 0;
disk_mem[ 3685] = 0;
disk_mem[ 3686] = 0;
disk_mem[ 3687] = 0;
disk_mem[ 3688] = 0;
disk_mem[ 3689] = 0;
disk_mem[ 3690] = 0;
disk_mem[ 3691] = 0;
disk_mem[ 3692] = 0;
disk_mem[ 3693] = 0;
disk_mem[ 3694] = 0;
disk_mem[ 3695] = 0;
disk_mem[ 3696] = 0;
disk_mem[ 3697] = 0;
disk_mem[ 3698] = 0;
disk_mem[ 3699] = 0;
disk_mem[ 3700] = 0;
disk_mem[ 3701] = 0;
disk_mem[ 3702] = 0;
disk_mem[ 3703] = 0;
disk_mem[ 3704] = 0;
disk_mem[ 3705] = 0;
disk_mem[ 3706] = 0;
disk_mem[ 3707] = 0;
disk_mem[ 3708] = 0;
disk_mem[ 3709] = 0;
disk_mem[ 3710] = 0;
disk_mem[ 3711] = 0;
disk_mem[ 3712] = 0;
disk_mem[ 3713] = 0;
disk_mem[ 3714] = 0;
disk_mem[ 3715] = 0;
disk_mem[ 3716] = 0;
disk_mem[ 3717] = 0;
disk_mem[ 3718] = 0;
disk_mem[ 3719] = 0;
disk_mem[ 3720] = 0;
disk_mem[ 3721] = 0;
disk_mem[ 3722] = 0;
disk_mem[ 3723] = 0;
disk_mem[ 3724] = 0;
disk_mem[ 3725] = 0;
disk_mem[ 3726] = 0;
disk_mem[ 3727] = 0;
disk_mem[ 3728] = 0;
disk_mem[ 3729] = 0;
disk_mem[ 3730] = 0;
disk_mem[ 3731] = 0;
disk_mem[ 3732] = 0;
disk_mem[ 3733] = 0;
disk_mem[ 3734] = 0;
disk_mem[ 3735] = 0;
disk_mem[ 3736] = 0;
disk_mem[ 3737] = 0;
disk_mem[ 3738] = 0;
disk_mem[ 3739] = 0;
disk_mem[ 3740] = 0;
disk_mem[ 3741] = 0;
disk_mem[ 3742] = 0;
disk_mem[ 3743] = 0;
disk_mem[ 3744] = 0;
disk_mem[ 3745] = 0;
disk_mem[ 3746] = 0;
disk_mem[ 3747] = 0;
disk_mem[ 3748] = 0;
disk_mem[ 3749] = 0;
disk_mem[ 3750] = 0;
disk_mem[ 3751] = 0;
disk_mem[ 3752] = 0;
disk_mem[ 3753] = 0;
disk_mem[ 3754] = 0;
disk_mem[ 3755] = 0;
disk_mem[ 3756] = 0;
disk_mem[ 3757] = 0;
disk_mem[ 3758] = 0;
disk_mem[ 3759] = 0;
disk_mem[ 3760] = 0;
disk_mem[ 3761] = 0;
disk_mem[ 3762] = 0;
disk_mem[ 3763] = 0;
disk_mem[ 3764] = 0;
disk_mem[ 3765] = 0;
disk_mem[ 3766] = 0;
disk_mem[ 3767] = 0;
disk_mem[ 3768] = 0;
disk_mem[ 3769] = 0;
disk_mem[ 3770] = 0;
disk_mem[ 3771] = 0;
disk_mem[ 3772] = 0;
disk_mem[ 3773] = 0;
disk_mem[ 3774] = 0;
disk_mem[ 3775] = 0;
disk_mem[ 3776] = 0;
disk_mem[ 3777] = 0;
disk_mem[ 3778] = 0;
disk_mem[ 3779] = 0;
disk_mem[ 3780] = 0;
disk_mem[ 3781] = 0;
disk_mem[ 3782] = 0;
disk_mem[ 3783] = 0;
disk_mem[ 3784] = 0;
disk_mem[ 3785] = 0;
disk_mem[ 3786] = 0;
disk_mem[ 3787] = 0;
disk_mem[ 3788] = 0;
disk_mem[ 3789] = 0;
disk_mem[ 3790] = 0;
disk_mem[ 3791] = 0;
disk_mem[ 3792] = 0;
disk_mem[ 3793] = 0;
disk_mem[ 3794] = 0;
disk_mem[ 3795] = 0;
disk_mem[ 3796] = 0;
disk_mem[ 3797] = 0;
disk_mem[ 3798] = 0;
disk_mem[ 3799] = 0;
disk_mem[ 3800] = 0;
disk_mem[ 3801] = 0;
disk_mem[ 3802] = 0;
disk_mem[ 3803] = 0;
disk_mem[ 3804] = 0;
disk_mem[ 3805] = 0;
disk_mem[ 3806] = 0;
disk_mem[ 3807] = 0;
disk_mem[ 3808] = 0;
disk_mem[ 3809] = 0;
disk_mem[ 3810] = 0;
disk_mem[ 3811] = 0;
disk_mem[ 3812] = 0;
disk_mem[ 3813] = 0;
disk_mem[ 3814] = 0;
disk_mem[ 3815] = 0;
disk_mem[ 3816] = 0;
disk_mem[ 3817] = 0;
disk_mem[ 3818] = 0;
disk_mem[ 3819] = 0;
disk_mem[ 3820] = 0;
disk_mem[ 3821] = 0;
disk_mem[ 3822] = 0;
disk_mem[ 3823] = 0;
disk_mem[ 3824] = 0;
disk_mem[ 3825] = 0;
disk_mem[ 3826] = 0;
disk_mem[ 3827] = 0;
disk_mem[ 3828] = 0;
disk_mem[ 3829] = 0;
disk_mem[ 3830] = 0;
disk_mem[ 3831] = 0;
disk_mem[ 3832] = 0;
disk_mem[ 3833] = 0;
disk_mem[ 3834] = 0;
disk_mem[ 3835] = 0;
disk_mem[ 3836] = 0;
disk_mem[ 3837] = 0;
disk_mem[ 3838] = 0;
disk_mem[ 3839] = 0;
disk_mem[ 3840] = 0;
disk_mem[ 3841] = 0;
disk_mem[ 3842] = 0;
disk_mem[ 3843] = 0;
disk_mem[ 3844] = 0;
disk_mem[ 3845] = 0;
disk_mem[ 3846] = 0;
disk_mem[ 3847] = 0;
disk_mem[ 3848] = 0;
disk_mem[ 3849] = 0;
disk_mem[ 3850] = 0;
disk_mem[ 3851] = 0;
disk_mem[ 3852] = 0;
disk_mem[ 3853] = 0;
disk_mem[ 3854] = 0;
disk_mem[ 3855] = 0;
disk_mem[ 3856] = 0;
disk_mem[ 3857] = 0;
disk_mem[ 3858] = 0;
disk_mem[ 3859] = 0;
disk_mem[ 3860] = 0;
disk_mem[ 3861] = 0;
disk_mem[ 3862] = 0;
disk_mem[ 3863] = 0;
disk_mem[ 3864] = 0;
disk_mem[ 3865] = 0;
disk_mem[ 3866] = 0;
disk_mem[ 3867] = 0;
disk_mem[ 3868] = 0;
disk_mem[ 3869] = 0;
disk_mem[ 3870] = 0;
disk_mem[ 3871] = 0;
disk_mem[ 3872] = 0;
disk_mem[ 3873] = 0;
disk_mem[ 3874] = 0;
disk_mem[ 3875] = 0;
disk_mem[ 3876] = 0;
disk_mem[ 3877] = 0;
disk_mem[ 3878] = 0;
disk_mem[ 3879] = 0;
disk_mem[ 3880] = 0;
disk_mem[ 3881] = 0;
disk_mem[ 3882] = 0;
disk_mem[ 3883] = 0;
disk_mem[ 3884] = 0;
disk_mem[ 3885] = 0;
disk_mem[ 3886] = 0;
disk_mem[ 3887] = 0;
disk_mem[ 3888] = 0;
disk_mem[ 3889] = 0;
disk_mem[ 3890] = 0;
disk_mem[ 3891] = 0;
disk_mem[ 3892] = 0;
disk_mem[ 3893] = 0;
disk_mem[ 3894] = 0;
disk_mem[ 3895] = 0;
disk_mem[ 3896] = 0;
disk_mem[ 3897] = 0;
disk_mem[ 3898] = 0;
disk_mem[ 3899] = 0;
disk_mem[ 3900] = 0;
disk_mem[ 3901] = 0;
disk_mem[ 3902] = 0;
disk_mem[ 3903] = 0;
disk_mem[ 3904] = 0;
disk_mem[ 3905] = 0;
disk_mem[ 3906] = 0;
disk_mem[ 3907] = 0;
disk_mem[ 3908] = 0;
disk_mem[ 3909] = 0;
disk_mem[ 3910] = 0;
disk_mem[ 3911] = 0;
disk_mem[ 3912] = 0;
disk_mem[ 3913] = 0;
disk_mem[ 3914] = 0;
disk_mem[ 3915] = 0;
disk_mem[ 3916] = 0;
disk_mem[ 3917] = 0;
disk_mem[ 3918] = 0;
disk_mem[ 3919] = 0;
disk_mem[ 3920] = 0;
disk_mem[ 3921] = 0;
disk_mem[ 3922] = 0;
disk_mem[ 3923] = 0;
disk_mem[ 3924] = 0;
disk_mem[ 3925] = 0;
disk_mem[ 3926] = 0;
disk_mem[ 3927] = 0;
disk_mem[ 3928] = 0;
disk_mem[ 3929] = 0;
disk_mem[ 3930] = 0;
disk_mem[ 3931] = 0;
disk_mem[ 3932] = 0;
disk_mem[ 3933] = 0;
disk_mem[ 3934] = 0;
disk_mem[ 3935] = 0;
disk_mem[ 3936] = 0;
disk_mem[ 3937] = 0;
disk_mem[ 3938] = 0;
disk_mem[ 3939] = 0;
disk_mem[ 3940] = 0;
disk_mem[ 3941] = 0;
disk_mem[ 3942] = 0;
disk_mem[ 3943] = 0;
disk_mem[ 3944] = 0;
disk_mem[ 3945] = 0;
disk_mem[ 3946] = 0;
disk_mem[ 3947] = 0;
disk_mem[ 3948] = 0;
disk_mem[ 3949] = 0;
disk_mem[ 3950] = 0;
disk_mem[ 3951] = 0;
disk_mem[ 3952] = 0;
disk_mem[ 3953] = 0;
disk_mem[ 3954] = 0;
disk_mem[ 3955] = 0;
disk_mem[ 3956] = 0;
disk_mem[ 3957] = 0;
disk_mem[ 3958] = 0;
disk_mem[ 3959] = 0;
disk_mem[ 3960] = 0;
disk_mem[ 3961] = 0;
disk_mem[ 3962] = 0;
disk_mem[ 3963] = 0;
disk_mem[ 3964] = 0;
disk_mem[ 3965] = 0;
disk_mem[ 3966] = 0;
disk_mem[ 3967] = 0;
disk_mem[ 3968] = 0;
disk_mem[ 3969] = 0;
disk_mem[ 3970] = 0;
disk_mem[ 3971] = 0;
disk_mem[ 3972] = 0;
disk_mem[ 3973] = 0;
disk_mem[ 3974] = 0;
disk_mem[ 3975] = 0;
disk_mem[ 3976] = 0;
disk_mem[ 3977] = 0;
disk_mem[ 3978] = 0;
disk_mem[ 3979] = 0;
disk_mem[ 3980] = 0;
disk_mem[ 3981] = 0;
disk_mem[ 3982] = 0;
disk_mem[ 3983] = 0;
disk_mem[ 3984] = 0;
disk_mem[ 3985] = 0;
disk_mem[ 3986] = 0;
disk_mem[ 3987] = 0;
disk_mem[ 3988] = 0;
disk_mem[ 3989] = 0;
disk_mem[ 3990] = 0;
disk_mem[ 3991] = 0;
disk_mem[ 3992] = 0;
disk_mem[ 3993] = 0;
disk_mem[ 3994] = 0;
disk_mem[ 3995] = 0;
disk_mem[ 3996] = 0;
disk_mem[ 3997] = 0;
disk_mem[ 3998] = 0;
disk_mem[ 3999] = 0;
disk_mem[ 4000] = 0;
disk_mem[ 4001] = 0;
disk_mem[ 4002] = 0;
disk_mem[ 4003] = 0;
disk_mem[ 4004] = 0;
disk_mem[ 4005] = 0;
disk_mem[ 4006] = 0;
disk_mem[ 4007] = 0;
disk_mem[ 4008] = 0;
disk_mem[ 4009] = 0;
disk_mem[ 4010] = 0;
disk_mem[ 4011] = 0;
disk_mem[ 4012] = 0;
disk_mem[ 4013] = 0;
disk_mem[ 4014] = 0;
disk_mem[ 4015] = 0;
disk_mem[ 4016] = 0;
disk_mem[ 4017] = 0;
disk_mem[ 4018] = 0;
disk_mem[ 4019] = 0;
disk_mem[ 4020] = 0;
disk_mem[ 4021] = 0;
disk_mem[ 4022] = 0;
disk_mem[ 4023] = 0;
disk_mem[ 4024] = 0;
disk_mem[ 4025] = 0;
disk_mem[ 4026] = 0;
disk_mem[ 4027] = 0;
disk_mem[ 4028] = 0;
disk_mem[ 4029] = 0;
disk_mem[ 4030] = 0;
disk_mem[ 4031] = 0;
disk_mem[ 4032] = 0;
disk_mem[ 4033] = 0;
disk_mem[ 4034] = 0;
disk_mem[ 4035] = 0;
disk_mem[ 4036] = 0;
disk_mem[ 4037] = 0;
disk_mem[ 4038] = 0;
disk_mem[ 4039] = 0;
disk_mem[ 4040] = 0;
disk_mem[ 4041] = 0;
disk_mem[ 4042] = 0;
disk_mem[ 4043] = 0;
disk_mem[ 4044] = 0;
disk_mem[ 4045] = 0;
disk_mem[ 4046] = 0;
disk_mem[ 4047] = 0;
disk_mem[ 4048] = 0;
disk_mem[ 4049] = 0;
disk_mem[ 4050] = 0;
disk_mem[ 4051] = 0;
disk_mem[ 4052] = 0;
disk_mem[ 4053] = 0;
disk_mem[ 4054] = 0;
disk_mem[ 4055] = 0;
disk_mem[ 4056] = 0;
disk_mem[ 4057] = 0;
disk_mem[ 4058] = 0;
disk_mem[ 4059] = 0;
disk_mem[ 4060] = 0;
disk_mem[ 4061] = 0;
disk_mem[ 4062] = 0;
disk_mem[ 4063] = 0;
disk_mem[ 4064] = 0;
disk_mem[ 4065] = 0;
disk_mem[ 4066] = 0;
disk_mem[ 4067] = 0;
disk_mem[ 4068] = 0;
disk_mem[ 4069] = 0;
disk_mem[ 4070] = 0;
disk_mem[ 4071] = 0;
disk_mem[ 4072] = 0;
disk_mem[ 4073] = 0;
disk_mem[ 4074] = 0;
disk_mem[ 4075] = 0;
disk_mem[ 4076] = 0;
disk_mem[ 4077] = 0;
disk_mem[ 4078] = 0;
disk_mem[ 4079] = 0;
disk_mem[ 4080] = 0;
disk_mem[ 4081] = 0;
disk_mem[ 4082] = 0;
disk_mem[ 4083] = 0;
disk_mem[ 4084] = 0;
disk_mem[ 4085] = 0;
disk_mem[ 4086] = 0;
disk_mem[ 4087] = 0;
disk_mem[ 4088] = 0;
disk_mem[ 4089] = 0;
disk_mem[ 4090] = 0;
disk_mem[ 4091] = 0;
disk_mem[ 4092] = 0;
disk_mem[ 4093] = 0;
disk_mem[ 4094] = 0;
disk_mem[ 4095] = 0;
disk_mem[ 4096] = 'hF8;
disk_mem[ 4097] = 'hFF;
disk_mem[ 4098] = 'hFF;
disk_mem[ 4099] = 'hFF;
disk_mem[ 4100] = 'hFF;
disk_mem[ 4101] = 'hFF;
disk_mem[ 4102] = 'hFF;
disk_mem[ 4103] = 'hFF;
disk_mem[ 4104] = 'hFF;
disk_mem[ 4105] = 0;
disk_mem[ 4106] = 0;
disk_mem[ 4107] = 0;
disk_mem[ 4108] = 0;
disk_mem[ 4109] = 0;
disk_mem[ 4110] = 0;
disk_mem[ 4111] = 0;
disk_mem[ 4112] = 0;
disk_mem[ 4113] = 0;
disk_mem[ 4114] = 0;
disk_mem[ 4115] = 0;
disk_mem[ 4116] = 0;
disk_mem[ 4117] = 0;
disk_mem[ 4118] = 0;
disk_mem[ 4119] = 0;
disk_mem[ 4120] = 0;
disk_mem[ 4121] = 0;
disk_mem[ 4122] = 0;
disk_mem[ 4123] = 0;
disk_mem[ 4124] = 0;
disk_mem[ 4125] = 0;
disk_mem[ 4126] = 0;
disk_mem[ 4127] = 0;
disk_mem[ 4128] = 0;
disk_mem[ 4129] = 0;
disk_mem[ 4130] = 0;
disk_mem[ 4131] = 0;
disk_mem[ 4132] = 0;
disk_mem[ 4133] = 0;
disk_mem[ 4134] = 0;
disk_mem[ 4135] = 0;
disk_mem[ 4136] = 0;
disk_mem[ 4137] = 0;
disk_mem[ 4138] = 0;
disk_mem[ 4139] = 0;
disk_mem[ 4140] = 0;
disk_mem[ 4141] = 0;
disk_mem[ 4142] = 0;
disk_mem[ 4143] = 0;
disk_mem[ 4144] = 0;
disk_mem[ 4145] = 0;
disk_mem[ 4146] = 0;
disk_mem[ 4147] = 0;
disk_mem[ 4148] = 0;
disk_mem[ 4149] = 0;
disk_mem[ 4150] = 0;
disk_mem[ 4151] = 0;
disk_mem[ 4152] = 0;
disk_mem[ 4153] = 0;
disk_mem[ 4154] = 0;
disk_mem[ 4155] = 0;
disk_mem[ 4156] = 0;
disk_mem[ 4157] = 0;
disk_mem[ 4158] = 0;
disk_mem[ 4159] = 0;
disk_mem[ 4160] = 0;
disk_mem[ 4161] = 0;
disk_mem[ 4162] = 0;
disk_mem[ 4163] = 0;
disk_mem[ 4164] = 0;
disk_mem[ 4165] = 0;
disk_mem[ 4166] = 0;
disk_mem[ 4167] = 0;
disk_mem[ 4168] = 0;
disk_mem[ 4169] = 0;
disk_mem[ 4170] = 0;
disk_mem[ 4171] = 0;
disk_mem[ 4172] = 0;
disk_mem[ 4173] = 0;
disk_mem[ 4174] = 0;
disk_mem[ 4175] = 0;
disk_mem[ 4176] = 0;
disk_mem[ 4177] = 0;
disk_mem[ 4178] = 0;
disk_mem[ 4179] = 0;
disk_mem[ 4180] = 0;
disk_mem[ 4181] = 0;
disk_mem[ 4182] = 0;
disk_mem[ 4183] = 0;
disk_mem[ 4184] = 0;
disk_mem[ 4185] = 0;
disk_mem[ 4186] = 0;
disk_mem[ 4187] = 0;
disk_mem[ 4188] = 0;
disk_mem[ 4189] = 0;
disk_mem[ 4190] = 0;
disk_mem[ 4191] = 0;
disk_mem[ 4192] = 0;
disk_mem[ 4193] = 0;
disk_mem[ 4194] = 0;
disk_mem[ 4195] = 0;
disk_mem[ 4196] = 0;
disk_mem[ 4197] = 0;
disk_mem[ 4198] = 0;
disk_mem[ 4199] = 0;
disk_mem[ 4200] = 0;
disk_mem[ 4201] = 0;
disk_mem[ 4202] = 0;
disk_mem[ 4203] = 0;
disk_mem[ 4204] = 0;
disk_mem[ 4205] = 0;
disk_mem[ 4206] = 0;
disk_mem[ 4207] = 0;
disk_mem[ 4208] = 0;
disk_mem[ 4209] = 0;
disk_mem[ 4210] = 0;
disk_mem[ 4211] = 0;
disk_mem[ 4212] = 0;
disk_mem[ 4213] = 0;
disk_mem[ 4214] = 0;
disk_mem[ 4215] = 0;
disk_mem[ 4216] = 0;
disk_mem[ 4217] = 0;
disk_mem[ 4218] = 0;
disk_mem[ 4219] = 0;
disk_mem[ 4220] = 0;
disk_mem[ 4221] = 0;
disk_mem[ 4222] = 0;
disk_mem[ 4223] = 0;
disk_mem[ 4224] = 0;
disk_mem[ 4225] = 0;
disk_mem[ 4226] = 0;
disk_mem[ 4227] = 0;
disk_mem[ 4228] = 0;
disk_mem[ 4229] = 0;
disk_mem[ 4230] = 0;
disk_mem[ 4231] = 0;
disk_mem[ 4232] = 0;
disk_mem[ 4233] = 0;
disk_mem[ 4234] = 0;
disk_mem[ 4235] = 0;
disk_mem[ 4236] = 0;
disk_mem[ 4237] = 0;
disk_mem[ 4238] = 0;
disk_mem[ 4239] = 0;
disk_mem[ 4240] = 0;
disk_mem[ 4241] = 0;
disk_mem[ 4242] = 0;
disk_mem[ 4243] = 0;
disk_mem[ 4244] = 0;
disk_mem[ 4245] = 0;
disk_mem[ 4246] = 0;
disk_mem[ 4247] = 0;
disk_mem[ 4248] = 0;
disk_mem[ 4249] = 0;
disk_mem[ 4250] = 0;
disk_mem[ 4251] = 0;
disk_mem[ 4252] = 0;
disk_mem[ 4253] = 0;
disk_mem[ 4254] = 0;
disk_mem[ 4255] = 0;
disk_mem[ 4256] = 0;
disk_mem[ 4257] = 0;
disk_mem[ 4258] = 0;
disk_mem[ 4259] = 0;
disk_mem[ 4260] = 0;
disk_mem[ 4261] = 0;
disk_mem[ 4262] = 0;
disk_mem[ 4263] = 0;
disk_mem[ 4264] = 0;
disk_mem[ 4265] = 0;
disk_mem[ 4266] = 0;
disk_mem[ 4267] = 0;
disk_mem[ 4268] = 0;
disk_mem[ 4269] = 0;
disk_mem[ 4270] = 0;
disk_mem[ 4271] = 0;
disk_mem[ 4272] = 0;
disk_mem[ 4273] = 0;
disk_mem[ 4274] = 0;
disk_mem[ 4275] = 0;
disk_mem[ 4276] = 0;
disk_mem[ 4277] = 0;
disk_mem[ 4278] = 0;
disk_mem[ 4279] = 0;
disk_mem[ 4280] = 0;
disk_mem[ 4281] = 0;
disk_mem[ 4282] = 0;
disk_mem[ 4283] = 0;
disk_mem[ 4284] = 0;
disk_mem[ 4285] = 0;
disk_mem[ 4286] = 0;
disk_mem[ 4287] = 0;
disk_mem[ 4288] = 0;
disk_mem[ 4289] = 0;
disk_mem[ 4290] = 0;
disk_mem[ 4291] = 0;
disk_mem[ 4292] = 0;
disk_mem[ 4293] = 0;
disk_mem[ 4294] = 0;
disk_mem[ 4295] = 0;
disk_mem[ 4296] = 0;
disk_mem[ 4297] = 0;
disk_mem[ 4298] = 0;
disk_mem[ 4299] = 0;
disk_mem[ 4300] = 0;
disk_mem[ 4301] = 0;
disk_mem[ 4302] = 0;
disk_mem[ 4303] = 0;
disk_mem[ 4304] = 0;
disk_mem[ 4305] = 0;
disk_mem[ 4306] = 0;
disk_mem[ 4307] = 0;
disk_mem[ 4308] = 0;
disk_mem[ 4309] = 0;
disk_mem[ 4310] = 0;
disk_mem[ 4311] = 0;
disk_mem[ 4312] = 0;
disk_mem[ 4313] = 0;
disk_mem[ 4314] = 0;
disk_mem[ 4315] = 0;
disk_mem[ 4316] = 0;
disk_mem[ 4317] = 0;
disk_mem[ 4318] = 0;
disk_mem[ 4319] = 0;
disk_mem[ 4320] = 0;
disk_mem[ 4321] = 0;
disk_mem[ 4322] = 0;
disk_mem[ 4323] = 0;
disk_mem[ 4324] = 0;
disk_mem[ 4325] = 0;
disk_mem[ 4326] = 0;
disk_mem[ 4327] = 0;
disk_mem[ 4328] = 0;
disk_mem[ 4329] = 0;
disk_mem[ 4330] = 0;
disk_mem[ 4331] = 0;
disk_mem[ 4332] = 0;
disk_mem[ 4333] = 0;
disk_mem[ 4334] = 0;
disk_mem[ 4335] = 0;
disk_mem[ 4336] = 0;
disk_mem[ 4337] = 0;
disk_mem[ 4338] = 0;
disk_mem[ 4339] = 0;
disk_mem[ 4340] = 0;
disk_mem[ 4341] = 0;
disk_mem[ 4342] = 0;
disk_mem[ 4343] = 0;
disk_mem[ 4344] = 0;
disk_mem[ 4345] = 0;
disk_mem[ 4346] = 0;
disk_mem[ 4347] = 0;
disk_mem[ 4348] = 0;
disk_mem[ 4349] = 0;
disk_mem[ 4350] = 0;
disk_mem[ 4351] = 0;
disk_mem[ 4352] = 0;
disk_mem[ 4353] = 0;
disk_mem[ 4354] = 0;
disk_mem[ 4355] = 0;
disk_mem[ 4356] = 0;
disk_mem[ 4357] = 0;
disk_mem[ 4358] = 0;
disk_mem[ 4359] = 0;
disk_mem[ 4360] = 0;
disk_mem[ 4361] = 0;
disk_mem[ 4362] = 0;
disk_mem[ 4363] = 0;
disk_mem[ 4364] = 0;
disk_mem[ 4365] = 0;
disk_mem[ 4366] = 0;
disk_mem[ 4367] = 0;
disk_mem[ 4368] = 0;
disk_mem[ 4369] = 0;
disk_mem[ 4370] = 0;
disk_mem[ 4371] = 0;
disk_mem[ 4372] = 0;
disk_mem[ 4373] = 0;
disk_mem[ 4374] = 0;
disk_mem[ 4375] = 0;
disk_mem[ 4376] = 0;
disk_mem[ 4377] = 0;
disk_mem[ 4378] = 0;
disk_mem[ 4379] = 0;
disk_mem[ 4380] = 0;
disk_mem[ 4381] = 0;
disk_mem[ 4382] = 0;
disk_mem[ 4383] = 0;
disk_mem[ 4384] = 0;
disk_mem[ 4385] = 0;
disk_mem[ 4386] = 0;
disk_mem[ 4387] = 0;
disk_mem[ 4388] = 0;
disk_mem[ 4389] = 0;
disk_mem[ 4390] = 0;
disk_mem[ 4391] = 0;
disk_mem[ 4392] = 0;
disk_mem[ 4393] = 0;
disk_mem[ 4394] = 0;
disk_mem[ 4395] = 0;
disk_mem[ 4396] = 0;
disk_mem[ 4397] = 0;
disk_mem[ 4398] = 0;
disk_mem[ 4399] = 0;
disk_mem[ 4400] = 0;
disk_mem[ 4401] = 0;
disk_mem[ 4402] = 0;
disk_mem[ 4403] = 0;
disk_mem[ 4404] = 0;
disk_mem[ 4405] = 0;
disk_mem[ 4406] = 0;
disk_mem[ 4407] = 0;
disk_mem[ 4408] = 0;
disk_mem[ 4409] = 0;
disk_mem[ 4410] = 0;
disk_mem[ 4411] = 0;
disk_mem[ 4412] = 0;
disk_mem[ 4413] = 0;
disk_mem[ 4414] = 0;
disk_mem[ 4415] = 0;
disk_mem[ 4416] = 0;
disk_mem[ 4417] = 0;
disk_mem[ 4418] = 0;
disk_mem[ 4419] = 0;
disk_mem[ 4420] = 0;
disk_mem[ 4421] = 0;
disk_mem[ 4422] = 0;
disk_mem[ 4423] = 0;
disk_mem[ 4424] = 0;
disk_mem[ 4425] = 0;
disk_mem[ 4426] = 0;
disk_mem[ 4427] = 0;
disk_mem[ 4428] = 0;
disk_mem[ 4429] = 0;
disk_mem[ 4430] = 0;
disk_mem[ 4431] = 0;
disk_mem[ 4432] = 0;
disk_mem[ 4433] = 0;
disk_mem[ 4434] = 0;
disk_mem[ 4435] = 0;
disk_mem[ 4436] = 0;
disk_mem[ 4437] = 0;
disk_mem[ 4438] = 0;
disk_mem[ 4439] = 0;
disk_mem[ 4440] = 0;
disk_mem[ 4441] = 0;
disk_mem[ 4442] = 0;
disk_mem[ 4443] = 0;
disk_mem[ 4444] = 0;
disk_mem[ 4445] = 0;
disk_mem[ 4446] = 0;
disk_mem[ 4447] = 0;
disk_mem[ 4448] = 0;
disk_mem[ 4449] = 0;
disk_mem[ 4450] = 0;
disk_mem[ 4451] = 0;
disk_mem[ 4452] = 0;
disk_mem[ 4453] = 0;
disk_mem[ 4454] = 0;
disk_mem[ 4455] = 0;
disk_mem[ 4456] = 0;
disk_mem[ 4457] = 0;
disk_mem[ 4458] = 0;
disk_mem[ 4459] = 0;
disk_mem[ 4460] = 0;
disk_mem[ 4461] = 0;
disk_mem[ 4462] = 0;
disk_mem[ 4463] = 0;
disk_mem[ 4464] = 0;
disk_mem[ 4465] = 0;
disk_mem[ 4466] = 0;
disk_mem[ 4467] = 0;
disk_mem[ 4468] = 0;
disk_mem[ 4469] = 0;
disk_mem[ 4470] = 0;
disk_mem[ 4471] = 0;
disk_mem[ 4472] = 0;
disk_mem[ 4473] = 0;
disk_mem[ 4474] = 0;
disk_mem[ 4475] = 0;
disk_mem[ 4476] = 0;
disk_mem[ 4477] = 0;
disk_mem[ 4478] = 0;
disk_mem[ 4479] = 0;
disk_mem[ 4480] = 0;
disk_mem[ 4481] = 0;
disk_mem[ 4482] = 0;
disk_mem[ 4483] = 0;
disk_mem[ 4484] = 0;
disk_mem[ 4485] = 0;
disk_mem[ 4486] = 0;
disk_mem[ 4487] = 0;
disk_mem[ 4488] = 0;
disk_mem[ 4489] = 0;
disk_mem[ 4490] = 0;
disk_mem[ 4491] = 0;
disk_mem[ 4492] = 0;
disk_mem[ 4493] = 0;
disk_mem[ 4494] = 0;
disk_mem[ 4495] = 0;
disk_mem[ 4496] = 0;
disk_mem[ 4497] = 0;
disk_mem[ 4498] = 0;
disk_mem[ 4499] = 0;
disk_mem[ 4500] = 0;
disk_mem[ 4501] = 0;
disk_mem[ 4502] = 0;
disk_mem[ 4503] = 0;
disk_mem[ 4504] = 0;
disk_mem[ 4505] = 0;
disk_mem[ 4506] = 0;
disk_mem[ 4507] = 0;
disk_mem[ 4508] = 0;
disk_mem[ 4509] = 0;
disk_mem[ 4510] = 0;
disk_mem[ 4511] = 0;
disk_mem[ 4512] = 0;
disk_mem[ 4513] = 0;
disk_mem[ 4514] = 0;
disk_mem[ 4515] = 0;
disk_mem[ 4516] = 0;
disk_mem[ 4517] = 0;
disk_mem[ 4518] = 0;
disk_mem[ 4519] = 0;
disk_mem[ 4520] = 0;
disk_mem[ 4521] = 0;
disk_mem[ 4522] = 0;
disk_mem[ 4523] = 0;
disk_mem[ 4524] = 0;
disk_mem[ 4525] = 0;
disk_mem[ 4526] = 0;
disk_mem[ 4527] = 0;
disk_mem[ 4528] = 0;
disk_mem[ 4529] = 0;
disk_mem[ 4530] = 0;
disk_mem[ 4531] = 0;
disk_mem[ 4532] = 0;
disk_mem[ 4533] = 0;
disk_mem[ 4534] = 0;
disk_mem[ 4535] = 0;
disk_mem[ 4536] = 0;
disk_mem[ 4537] = 0;
disk_mem[ 4538] = 0;
disk_mem[ 4539] = 0;
disk_mem[ 4540] = 0;
disk_mem[ 4541] = 0;
disk_mem[ 4542] = 0;
disk_mem[ 4543] = 0;
disk_mem[ 4544] = 0;
disk_mem[ 4545] = 0;
disk_mem[ 4546] = 0;
disk_mem[ 4547] = 0;
disk_mem[ 4548] = 0;
disk_mem[ 4549] = 0;
disk_mem[ 4550] = 0;
disk_mem[ 4551] = 0;
disk_mem[ 4552] = 0;
disk_mem[ 4553] = 0;
disk_mem[ 4554] = 0;
disk_mem[ 4555] = 0;
disk_mem[ 4556] = 0;
disk_mem[ 4557] = 0;
disk_mem[ 4558] = 0;
disk_mem[ 4559] = 0;
disk_mem[ 4560] = 0;
disk_mem[ 4561] = 0;
disk_mem[ 4562] = 0;
disk_mem[ 4563] = 0;
disk_mem[ 4564] = 0;
disk_mem[ 4565] = 0;
disk_mem[ 4566] = 0;
disk_mem[ 4567] = 0;
disk_mem[ 4568] = 0;
disk_mem[ 4569] = 0;
disk_mem[ 4570] = 0;
disk_mem[ 4571] = 0;
disk_mem[ 4572] = 0;
disk_mem[ 4573] = 0;
disk_mem[ 4574] = 0;
disk_mem[ 4575] = 0;
disk_mem[ 4576] = 0;
disk_mem[ 4577] = 0;
disk_mem[ 4578] = 0;
disk_mem[ 4579] = 0;
disk_mem[ 4580] = 0;
disk_mem[ 4581] = 0;
disk_mem[ 4582] = 0;
disk_mem[ 4583] = 0;
disk_mem[ 4584] = 0;
disk_mem[ 4585] = 0;
disk_mem[ 4586] = 0;
disk_mem[ 4587] = 0;
disk_mem[ 4588] = 0;
disk_mem[ 4589] = 0;
disk_mem[ 4590] = 0;
disk_mem[ 4591] = 0;
disk_mem[ 4592] = 0;
disk_mem[ 4593] = 0;
disk_mem[ 4594] = 0;
disk_mem[ 4595] = 0;
disk_mem[ 4596] = 0;
disk_mem[ 4597] = 0;
disk_mem[ 4598] = 0;
disk_mem[ 4599] = 0;
disk_mem[ 4600] = 0;
disk_mem[ 4601] = 0;
disk_mem[ 4602] = 0;
disk_mem[ 4603] = 0;
disk_mem[ 4604] = 0;
disk_mem[ 4605] = 0;
disk_mem[ 4606] = 0;
disk_mem[ 4607] = 0;
disk_mem[ 4608] = 'h42;
disk_mem[ 4609] = 'h20;
disk_mem[ 4610] = 0;
disk_mem[ 4611] = 'h49;
disk_mem[ 4612] = 0;
disk_mem[ 4613] = 'h6E;
disk_mem[ 4614] = 0;
disk_mem[ 4615] = 'h66;
disk_mem[ 4616] = 0;
disk_mem[ 4617] = 'h6F;
disk_mem[ 4618] = 0;
disk_mem[ 4619] = 'h0F;
disk_mem[ 4620] = 0;
disk_mem[ 4621] = 'h72;
disk_mem[ 4622] = 'h72;
disk_mem[ 4623] = 0;
disk_mem[ 4624] = 'h6D;
disk_mem[ 4625] = 0;
disk_mem[ 4626] = 'h61;
disk_mem[ 4627] = 0;
disk_mem[ 4628] = 'h74;
disk_mem[ 4629] = 0;
disk_mem[ 4630] = 'h69;
disk_mem[ 4631] = 0;
disk_mem[ 4632] = 'h6F;
disk_mem[ 4633] = 0;
disk_mem[ 4634] = 0;
disk_mem[ 4635] = 0;
disk_mem[ 4636] = 'h6E;
disk_mem[ 4637] = 0;
disk_mem[ 4638] = 0;
disk_mem[ 4639] = 0;
disk_mem[ 4640] = 'h01;
disk_mem[ 4641] = 'h53;
disk_mem[ 4642] = 0;
disk_mem[ 4643] = 'h79;
disk_mem[ 4644] = 0;
disk_mem[ 4645] = 'h73;
disk_mem[ 4646] = 0;
disk_mem[ 4647] = 'h74;
disk_mem[ 4648] = 0;
disk_mem[ 4649] = 'h65;
disk_mem[ 4650] = 0;
disk_mem[ 4651] = 'h0F;
disk_mem[ 4652] = 0;
disk_mem[ 4653] = 'h72;
disk_mem[ 4654] = 'h6D;
disk_mem[ 4655] = 0;
disk_mem[ 4656] = 'h20;
disk_mem[ 4657] = 0;
disk_mem[ 4658] = 'h56;
disk_mem[ 4659] = 0;
disk_mem[ 4660] = 'h6F;
disk_mem[ 4661] = 0;
disk_mem[ 4662] = 'h6C;
disk_mem[ 4663] = 0;
disk_mem[ 4664] = 'h75;
disk_mem[ 4665] = 0;
disk_mem[ 4666] = 0;
disk_mem[ 4667] = 0;
disk_mem[ 4668] = 'h6D;
disk_mem[ 4669] = 0;
disk_mem[ 4670] = 'h65;
disk_mem[ 4671] = 0;
disk_mem[ 4672] = 'h53;
disk_mem[ 4673] = 'h59;
disk_mem[ 4674] = 'h53;
disk_mem[ 4675] = 'h54;
disk_mem[ 4676] = 'h45;
disk_mem[ 4677] = 'h4D;
disk_mem[ 4678] = 'h7E;
disk_mem[ 4679] = 'h31;
disk_mem[ 4680] = 'h20;
disk_mem[ 4681] = 'h20;
disk_mem[ 4682] = 'h20;
disk_mem[ 4683] = 'h16;
disk_mem[ 4684] = 0;
disk_mem[ 4685] = 'h8B;
disk_mem[ 4686] = 'h90;
disk_mem[ 4687] = 'h80;
disk_mem[ 4688] = 'h43;
disk_mem[ 4689] = 'h55;
disk_mem[ 4690] = 'h43;
disk_mem[ 4691] = 'h55;
disk_mem[ 4692] = 0;
disk_mem[ 4693] = 0;
disk_mem[ 4694] = 'h91;
disk_mem[ 4695] = 'h80;
disk_mem[ 4696] = 'h43;
disk_mem[ 4697] = 'h55;
disk_mem[ 4698] = 'h02;
disk_mem[ 4699] = 0;
disk_mem[ 4700] = 0;
disk_mem[ 4701] = 0;
disk_mem[ 4702] = 0;
disk_mem[ 4703] = 0;
disk_mem[ 4704] = 'h45;
disk_mem[ 4705] = 'h58;
disk_mem[ 4706] = 'h41;
disk_mem[ 4707] = 'h4D;
disk_mem[ 4708] = 'h50;
disk_mem[ 4709] = 'h4C;
disk_mem[ 4710] = 'h45;
disk_mem[ 4711] = 'h20;
disk_mem[ 4712] = 'h54;
disk_mem[ 4713] = 'h58;
disk_mem[ 4714] = 'h54;
disk_mem[ 4715] = 'h20;
disk_mem[ 4716] = 'h18;
disk_mem[ 4717] = 'h1C;
disk_mem[ 4718] = 'h9A;
disk_mem[ 4719] = 'h80;
disk_mem[ 4720] = 'h43;
disk_mem[ 4721] = 'h55;
disk_mem[ 4722] = 'h43;
disk_mem[ 4723] = 'h55;
disk_mem[ 4724] = 0;
disk_mem[ 4725] = 0;
disk_mem[ 4726] = 'hAF;
disk_mem[ 4727] = 'h80;
disk_mem[ 4728] = 'h43;
disk_mem[ 4729] = 'h55;
disk_mem[ 4730] = 'h05;
disk_mem[ 4731] = 0;
disk_mem[ 4732] = 'h26;
disk_mem[ 4733] = 0;
disk_mem[ 4734] = 0;
disk_mem[ 4735] = 0;
disk_mem[ 4736] = 0;
disk_mem[ 4737] = 0;
disk_mem[ 4738] = 0;
disk_mem[ 4739] = 0;
disk_mem[ 4740] = 0;
disk_mem[ 4741] = 0;
disk_mem[ 4742] = 0;
disk_mem[ 4743] = 0;
disk_mem[ 4744] = 0;
disk_mem[ 4745] = 0;
disk_mem[ 4746] = 0;
disk_mem[ 4747] = 0;
disk_mem[ 4748] = 0;
disk_mem[ 4749] = 0;
disk_mem[ 4750] = 0;
disk_mem[ 4751] = 0;
disk_mem[ 4752] = 0;
disk_mem[ 4753] = 0;
disk_mem[ 4754] = 0;
disk_mem[ 4755] = 0;
disk_mem[ 4756] = 0;
disk_mem[ 4757] = 0;
disk_mem[ 4758] = 0;
disk_mem[ 4759] = 0;
disk_mem[ 4760] = 0;
disk_mem[ 4761] = 0;
disk_mem[ 4762] = 0;
disk_mem[ 4763] = 0;
disk_mem[ 4764] = 0;
disk_mem[ 4765] = 0;
disk_mem[ 4766] = 0;
disk_mem[ 4767] = 0;
disk_mem[ 4768] = 0;
disk_mem[ 4769] = 0;
disk_mem[ 4770] = 0;
disk_mem[ 4771] = 0;
disk_mem[ 4772] = 0;
disk_mem[ 4773] = 0;
disk_mem[ 4774] = 0;
disk_mem[ 4775] = 0;
disk_mem[ 4776] = 0;
disk_mem[ 4777] = 0;
disk_mem[ 4778] = 0;
disk_mem[ 4779] = 0;
disk_mem[ 4780] = 0;
disk_mem[ 4781] = 0;
disk_mem[ 4782] = 0;
disk_mem[ 4783] = 0;
disk_mem[ 4784] = 0;
disk_mem[ 4785] = 0;
disk_mem[ 4786] = 0;
disk_mem[ 4787] = 0;
disk_mem[ 4788] = 0;
disk_mem[ 4789] = 0;
disk_mem[ 4790] = 0;
disk_mem[ 4791] = 0;
disk_mem[ 4792] = 0;
disk_mem[ 4793] = 0;
disk_mem[ 4794] = 0;
disk_mem[ 4795] = 0;
disk_mem[ 4796] = 0;
disk_mem[ 4797] = 0;
disk_mem[ 4798] = 0;
disk_mem[ 4799] = 0;
disk_mem[ 4800] = 0;
disk_mem[ 4801] = 0;
disk_mem[ 4802] = 0;
disk_mem[ 4803] = 0;
disk_mem[ 4804] = 0;
disk_mem[ 4805] = 0;
disk_mem[ 4806] = 0;
disk_mem[ 4807] = 0;
disk_mem[ 4808] = 0;
disk_mem[ 4809] = 0;
disk_mem[ 4810] = 0;
disk_mem[ 4811] = 0;
disk_mem[ 4812] = 0;
disk_mem[ 4813] = 0;
disk_mem[ 4814] = 0;
disk_mem[ 4815] = 0;
disk_mem[ 4816] = 0;
disk_mem[ 4817] = 0;
disk_mem[ 4818] = 0;
disk_mem[ 4819] = 0;
disk_mem[ 4820] = 0;
disk_mem[ 4821] = 0;
disk_mem[ 4822] = 0;
disk_mem[ 4823] = 0;
disk_mem[ 4824] = 0;
disk_mem[ 4825] = 0;
disk_mem[ 4826] = 0;
disk_mem[ 4827] = 0;
disk_mem[ 4828] = 0;
disk_mem[ 4829] = 0;
disk_mem[ 4830] = 0;
disk_mem[ 4831] = 0;
disk_mem[ 4832] = 0;
disk_mem[ 4833] = 0;
disk_mem[ 4834] = 0;
disk_mem[ 4835] = 0;
disk_mem[ 4836] = 0;
disk_mem[ 4837] = 0;
disk_mem[ 4838] = 0;
disk_mem[ 4839] = 0;
disk_mem[ 4840] = 0;
disk_mem[ 4841] = 0;
disk_mem[ 4842] = 0;
disk_mem[ 4843] = 0;
disk_mem[ 4844] = 0;
disk_mem[ 4845] = 0;
disk_mem[ 4846] = 0;
disk_mem[ 4847] = 0;
disk_mem[ 4848] = 0;
disk_mem[ 4849] = 0;
disk_mem[ 4850] = 0;
disk_mem[ 4851] = 0;
disk_mem[ 4852] = 0;
disk_mem[ 4853] = 0;
disk_mem[ 4854] = 0;
disk_mem[ 4855] = 0;
disk_mem[ 4856] = 0;
disk_mem[ 4857] = 0;
disk_mem[ 4858] = 0;
disk_mem[ 4859] = 0;
disk_mem[ 4860] = 0;
disk_mem[ 4861] = 0;
disk_mem[ 4862] = 0;
disk_mem[ 4863] = 0;
disk_mem[ 4864] = 0;
disk_mem[ 4865] = 0;
disk_mem[ 4866] = 0;
disk_mem[ 4867] = 0;
disk_mem[ 4868] = 0;
disk_mem[ 4869] = 0;
disk_mem[ 4870] = 0;
disk_mem[ 4871] = 0;
disk_mem[ 4872] = 0;
disk_mem[ 4873] = 0;
disk_mem[ 4874] = 0;
disk_mem[ 4875] = 0;
disk_mem[ 4876] = 0;
disk_mem[ 4877] = 0;
disk_mem[ 4878] = 0;
disk_mem[ 4879] = 0;
disk_mem[ 4880] = 0;
disk_mem[ 4881] = 0;
disk_mem[ 4882] = 0;
disk_mem[ 4883] = 0;
disk_mem[ 4884] = 0;
disk_mem[ 4885] = 0;
disk_mem[ 4886] = 0;
disk_mem[ 4887] = 0;
disk_mem[ 4888] = 0;
disk_mem[ 4889] = 0;
disk_mem[ 4890] = 0;
disk_mem[ 4891] = 0;
disk_mem[ 4892] = 0;
disk_mem[ 4893] = 0;
disk_mem[ 4894] = 0;
disk_mem[ 4895] = 0;
disk_mem[ 4896] = 0;
disk_mem[ 4897] = 0;
disk_mem[ 4898] = 0;
disk_mem[ 4899] = 0;
disk_mem[ 4900] = 0;
disk_mem[ 4901] = 0;
disk_mem[ 4902] = 0;
disk_mem[ 4903] = 0;
disk_mem[ 4904] = 0;
disk_mem[ 4905] = 0;
disk_mem[ 4906] = 0;
disk_mem[ 4907] = 0;
disk_mem[ 4908] = 0;
disk_mem[ 4909] = 0;
disk_mem[ 4910] = 0;
disk_mem[ 4911] = 0;
disk_mem[ 4912] = 0;
disk_mem[ 4913] = 0;
disk_mem[ 4914] = 0;
disk_mem[ 4915] = 0;
disk_mem[ 4916] = 0;
disk_mem[ 4917] = 0;
disk_mem[ 4918] = 0;
disk_mem[ 4919] = 0;
disk_mem[ 4920] = 0;
disk_mem[ 4921] = 0;
disk_mem[ 4922] = 0;
disk_mem[ 4923] = 0;
disk_mem[ 4924] = 0;
disk_mem[ 4925] = 0;
disk_mem[ 4926] = 0;
disk_mem[ 4927] = 0;
disk_mem[ 4928] = 0;
disk_mem[ 4929] = 0;
disk_mem[ 4930] = 0;
disk_mem[ 4931] = 0;
disk_mem[ 4932] = 0;
disk_mem[ 4933] = 0;
disk_mem[ 4934] = 0;
disk_mem[ 4935] = 0;
disk_mem[ 4936] = 0;
disk_mem[ 4937] = 0;
disk_mem[ 4938] = 0;
disk_mem[ 4939] = 0;
disk_mem[ 4940] = 0;
disk_mem[ 4941] = 0;
disk_mem[ 4942] = 0;
disk_mem[ 4943] = 0;
disk_mem[ 4944] = 0;
disk_mem[ 4945] = 0;
disk_mem[ 4946] = 0;
disk_mem[ 4947] = 0;
disk_mem[ 4948] = 0;
disk_mem[ 4949] = 0;
disk_mem[ 4950] = 0;
disk_mem[ 4951] = 0;
disk_mem[ 4952] = 0;
disk_mem[ 4953] = 0;
disk_mem[ 4954] = 0;
disk_mem[ 4955] = 0;
disk_mem[ 4956] = 0;
disk_mem[ 4957] = 0;
disk_mem[ 4958] = 0;
disk_mem[ 4959] = 0;
disk_mem[ 4960] = 0;
disk_mem[ 4961] = 0;
disk_mem[ 4962] = 0;
disk_mem[ 4963] = 0;
disk_mem[ 4964] = 0;
disk_mem[ 4965] = 0;
disk_mem[ 4966] = 0;
disk_mem[ 4967] = 0;
disk_mem[ 4968] = 0;
disk_mem[ 4969] = 0;
disk_mem[ 4970] = 0;
disk_mem[ 4971] = 0;
disk_mem[ 4972] = 0;
disk_mem[ 4973] = 0;
disk_mem[ 4974] = 0;
disk_mem[ 4975] = 0;
disk_mem[ 4976] = 0;
disk_mem[ 4977] = 0;
disk_mem[ 4978] = 0;
disk_mem[ 4979] = 0;
disk_mem[ 4980] = 0;
disk_mem[ 4981] = 0;
disk_mem[ 4982] = 0;
disk_mem[ 4983] = 0;
disk_mem[ 4984] = 0;
disk_mem[ 4985] = 0;
disk_mem[ 4986] = 0;
disk_mem[ 4987] = 0;
disk_mem[ 4988] = 0;
disk_mem[ 4989] = 0;
disk_mem[ 4990] = 0;
disk_mem[ 4991] = 0;
disk_mem[ 4992] = 0;
disk_mem[ 4993] = 0;
disk_mem[ 4994] = 0;
disk_mem[ 4995] = 0;
disk_mem[ 4996] = 0;
disk_mem[ 4997] = 0;
disk_mem[ 4998] = 0;
disk_mem[ 4999] = 0;
disk_mem[ 5000] = 0;
disk_mem[ 5001] = 0;
disk_mem[ 5002] = 0;
disk_mem[ 5003] = 0;
disk_mem[ 5004] = 0;
disk_mem[ 5005] = 0;
disk_mem[ 5006] = 0;
disk_mem[ 5007] = 0;
disk_mem[ 5008] = 0;
disk_mem[ 5009] = 0;
disk_mem[ 5010] = 0;
disk_mem[ 5011] = 0;
disk_mem[ 5012] = 0;
disk_mem[ 5013] = 0;
disk_mem[ 5014] = 0;
disk_mem[ 5015] = 0;
disk_mem[ 5016] = 0;
disk_mem[ 5017] = 0;
disk_mem[ 5018] = 0;
disk_mem[ 5019] = 0;
disk_mem[ 5020] = 0;
disk_mem[ 5021] = 0;
disk_mem[ 5022] = 0;
disk_mem[ 5023] = 0;
disk_mem[ 5024] = 0;
disk_mem[ 5025] = 0;
disk_mem[ 5026] = 0;
disk_mem[ 5027] = 0;
disk_mem[ 5028] = 0;
disk_mem[ 5029] = 0;
disk_mem[ 5030] = 0;
disk_mem[ 5031] = 0;
disk_mem[ 5032] = 0;
disk_mem[ 5033] = 0;
disk_mem[ 5034] = 0;
disk_mem[ 5035] = 0;
disk_mem[ 5036] = 0;
disk_mem[ 5037] = 0;
disk_mem[ 5038] = 0;
disk_mem[ 5039] = 0;
disk_mem[ 5040] = 0;
disk_mem[ 5041] = 0;
disk_mem[ 5042] = 0;
disk_mem[ 5043] = 0;
disk_mem[ 5044] = 0;
disk_mem[ 5045] = 0;
disk_mem[ 5046] = 0;
disk_mem[ 5047] = 0;
disk_mem[ 5048] = 0;
disk_mem[ 5049] = 0;
disk_mem[ 5050] = 0;
disk_mem[ 5051] = 0;
disk_mem[ 5052] = 0;
disk_mem[ 5053] = 0;
disk_mem[ 5054] = 0;
disk_mem[ 5055] = 0;
disk_mem[ 5056] = 0;
disk_mem[ 5057] = 0;
disk_mem[ 5058] = 0;
disk_mem[ 5059] = 0;
disk_mem[ 5060] = 0;
disk_mem[ 5061] = 0;
disk_mem[ 5062] = 0;
disk_mem[ 5063] = 0;
disk_mem[ 5064] = 0;
disk_mem[ 5065] = 0;
disk_mem[ 5066] = 0;
disk_mem[ 5067] = 0;
disk_mem[ 5068] = 0;
disk_mem[ 5069] = 0;
disk_mem[ 5070] = 0;
disk_mem[ 5071] = 0;
disk_mem[ 5072] = 0;
disk_mem[ 5073] = 0;
disk_mem[ 5074] = 0;
disk_mem[ 5075] = 0;
disk_mem[ 5076] = 0;
disk_mem[ 5077] = 0;
disk_mem[ 5078] = 0;
disk_mem[ 5079] = 0;
disk_mem[ 5080] = 0;
disk_mem[ 5081] = 0;
disk_mem[ 5082] = 0;
disk_mem[ 5083] = 0;
disk_mem[ 5084] = 0;
disk_mem[ 5085] = 0;
disk_mem[ 5086] = 0;
disk_mem[ 5087] = 0;
disk_mem[ 5088] = 0;
disk_mem[ 5089] = 0;
disk_mem[ 5090] = 0;
disk_mem[ 5091] = 0;
disk_mem[ 5092] = 0;
disk_mem[ 5093] = 0;
disk_mem[ 5094] = 0;
disk_mem[ 5095] = 0;
disk_mem[ 5096] = 0;
disk_mem[ 5097] = 0;
disk_mem[ 5098] = 0;
disk_mem[ 5099] = 0;
disk_mem[ 5100] = 0;
disk_mem[ 5101] = 0;
disk_mem[ 5102] = 0;
disk_mem[ 5103] = 0;
disk_mem[ 5104] = 0;
disk_mem[ 5105] = 0;
disk_mem[ 5106] = 0;
disk_mem[ 5107] = 0;
disk_mem[ 5108] = 0;
disk_mem[ 5109] = 0;
disk_mem[ 5110] = 0;
disk_mem[ 5111] = 0;
disk_mem[ 5112] = 0;
disk_mem[ 5113] = 0;
disk_mem[ 5114] = 0;
disk_mem[ 5115] = 0;
disk_mem[ 5116] = 0;
disk_mem[ 5117] = 0;
disk_mem[ 5118] = 0;
disk_mem[ 5119] = 0;
disk_mem[ 5120] = 0;
disk_mem[ 5121] = 0;
disk_mem[ 5122] = 0;
disk_mem[ 5123] = 0;
disk_mem[ 5124] = 0;
disk_mem[ 5125] = 0;
disk_mem[ 5126] = 0;
disk_mem[ 5127] = 0;
disk_mem[ 5128] = 0;
disk_mem[ 5129] = 0;
disk_mem[ 5130] = 0;
disk_mem[ 5131] = 0;
disk_mem[ 5132] = 0;
disk_mem[ 5133] = 0;
disk_mem[ 5134] = 0;
disk_mem[ 5135] = 0;
disk_mem[ 5136] = 0;
disk_mem[ 5137] = 0;
disk_mem[ 5138] = 0;
disk_mem[ 5139] = 0;
disk_mem[ 5140] = 0;
disk_mem[ 5141] = 0;
disk_mem[ 5142] = 0;
disk_mem[ 5143] = 0;
disk_mem[ 5144] = 0;
disk_mem[ 5145] = 0;
disk_mem[ 5146] = 0;
disk_mem[ 5147] = 0;
disk_mem[ 5148] = 0;
disk_mem[ 5149] = 0;
disk_mem[ 5150] = 0;
disk_mem[ 5151] = 0;
disk_mem[ 5152] = 0;
disk_mem[ 5153] = 0;
disk_mem[ 5154] = 0;
disk_mem[ 5155] = 0;
disk_mem[ 5156] = 0;
disk_mem[ 5157] = 0;
disk_mem[ 5158] = 0;
disk_mem[ 5159] = 0;
disk_mem[ 5160] = 0;
disk_mem[ 5161] = 0;
disk_mem[ 5162] = 0;
disk_mem[ 5163] = 0;
disk_mem[ 5164] = 0;
disk_mem[ 5165] = 0;
disk_mem[ 5166] = 0;
disk_mem[ 5167] = 0;
disk_mem[ 5168] = 0;
disk_mem[ 5169] = 0;
disk_mem[ 5170] = 0;
disk_mem[ 5171] = 0;
disk_mem[ 5172] = 0;
disk_mem[ 5173] = 0;
disk_mem[ 5174] = 0;
disk_mem[ 5175] = 0;
disk_mem[ 5176] = 0;
disk_mem[ 5177] = 0;
disk_mem[ 5178] = 0;
disk_mem[ 5179] = 0;
disk_mem[ 5180] = 0;
disk_mem[ 5181] = 0;
disk_mem[ 5182] = 0;
disk_mem[ 5183] = 0;
disk_mem[ 5184] = 0;
disk_mem[ 5185] = 0;
disk_mem[ 5186] = 0;
disk_mem[ 5187] = 0;
disk_mem[ 5188] = 0;
disk_mem[ 5189] = 0;
disk_mem[ 5190] = 0;
disk_mem[ 5191] = 0;
disk_mem[ 5192] = 0;
disk_mem[ 5193] = 0;
disk_mem[ 5194] = 0;
disk_mem[ 5195] = 0;
disk_mem[ 5196] = 0;
disk_mem[ 5197] = 0;
disk_mem[ 5198] = 0;
disk_mem[ 5199] = 0;
disk_mem[ 5200] = 0;
disk_mem[ 5201] = 0;
disk_mem[ 5202] = 0;
disk_mem[ 5203] = 0;
disk_mem[ 5204] = 0;
disk_mem[ 5205] = 0;
disk_mem[ 5206] = 0;
disk_mem[ 5207] = 0;
disk_mem[ 5208] = 0;
disk_mem[ 5209] = 0;
disk_mem[ 5210] = 0;
disk_mem[ 5211] = 0;
disk_mem[ 5212] = 0;
disk_mem[ 5213] = 0;
disk_mem[ 5214] = 0;
disk_mem[ 5215] = 0;
disk_mem[ 5216] = 0;
disk_mem[ 5217] = 0;
disk_mem[ 5218] = 0;
disk_mem[ 5219] = 0;
disk_mem[ 5220] = 0;
disk_mem[ 5221] = 0;
disk_mem[ 5222] = 0;
disk_mem[ 5223] = 0;
disk_mem[ 5224] = 0;
disk_mem[ 5225] = 0;
disk_mem[ 5226] = 0;
disk_mem[ 5227] = 0;
disk_mem[ 5228] = 0;
disk_mem[ 5229] = 0;
disk_mem[ 5230] = 0;
disk_mem[ 5231] = 0;
disk_mem[ 5232] = 0;
disk_mem[ 5233] = 0;
disk_mem[ 5234] = 0;
disk_mem[ 5235] = 0;
disk_mem[ 5236] = 0;
disk_mem[ 5237] = 0;
disk_mem[ 5238] = 0;
disk_mem[ 5239] = 0;
disk_mem[ 5240] = 0;
disk_mem[ 5241] = 0;
disk_mem[ 5242] = 0;
disk_mem[ 5243] = 0;
disk_mem[ 5244] = 0;
disk_mem[ 5245] = 0;
disk_mem[ 5246] = 0;
disk_mem[ 5247] = 0;
disk_mem[ 5248] = 0;
disk_mem[ 5249] = 0;
disk_mem[ 5250] = 0;
disk_mem[ 5251] = 0;
disk_mem[ 5252] = 0;
disk_mem[ 5253] = 0;
disk_mem[ 5254] = 0;
disk_mem[ 5255] = 0;
disk_mem[ 5256] = 0;
disk_mem[ 5257] = 0;
disk_mem[ 5258] = 0;
disk_mem[ 5259] = 0;
disk_mem[ 5260] = 0;
disk_mem[ 5261] = 0;
disk_mem[ 5262] = 0;
disk_mem[ 5263] = 0;
disk_mem[ 5264] = 0;
disk_mem[ 5265] = 0;
disk_mem[ 5266] = 0;
disk_mem[ 5267] = 0;
disk_mem[ 5268] = 0;
disk_mem[ 5269] = 0;
disk_mem[ 5270] = 0;
disk_mem[ 5271] = 0;
disk_mem[ 5272] = 0;
disk_mem[ 5273] = 0;
disk_mem[ 5274] = 0;
disk_mem[ 5275] = 0;
disk_mem[ 5276] = 0;
disk_mem[ 5277] = 0;
disk_mem[ 5278] = 0;
disk_mem[ 5279] = 0;
disk_mem[ 5280] = 0;
disk_mem[ 5281] = 0;
disk_mem[ 5282] = 0;
disk_mem[ 5283] = 0;
disk_mem[ 5284] = 0;
disk_mem[ 5285] = 0;
disk_mem[ 5286] = 0;
disk_mem[ 5287] = 0;
disk_mem[ 5288] = 0;
disk_mem[ 5289] = 0;
disk_mem[ 5290] = 0;
disk_mem[ 5291] = 0;
disk_mem[ 5292] = 0;
disk_mem[ 5293] = 0;
disk_mem[ 5294] = 0;
disk_mem[ 5295] = 0;
disk_mem[ 5296] = 0;
disk_mem[ 5297] = 0;
disk_mem[ 5298] = 0;
disk_mem[ 5299] = 0;
disk_mem[ 5300] = 0;
disk_mem[ 5301] = 0;
disk_mem[ 5302] = 0;
disk_mem[ 5303] = 0;
disk_mem[ 5304] = 0;
disk_mem[ 5305] = 0;
disk_mem[ 5306] = 0;
disk_mem[ 5307] = 0;
disk_mem[ 5308] = 0;
disk_mem[ 5309] = 0;
disk_mem[ 5310] = 0;
disk_mem[ 5311] = 0;
disk_mem[ 5312] = 0;
disk_mem[ 5313] = 0;
disk_mem[ 5314] = 0;
disk_mem[ 5315] = 0;
disk_mem[ 5316] = 0;
disk_mem[ 5317] = 0;
disk_mem[ 5318] = 0;
disk_mem[ 5319] = 0;
disk_mem[ 5320] = 0;
disk_mem[ 5321] = 0;
disk_mem[ 5322] = 0;
disk_mem[ 5323] = 0;
disk_mem[ 5324] = 0;
disk_mem[ 5325] = 0;
disk_mem[ 5326] = 0;
disk_mem[ 5327] = 0;
disk_mem[ 5328] = 0;
disk_mem[ 5329] = 0;
disk_mem[ 5330] = 0;
disk_mem[ 5331] = 0;
disk_mem[ 5332] = 0;
disk_mem[ 5333] = 0;
disk_mem[ 5334] = 0;
disk_mem[ 5335] = 0;
disk_mem[ 5336] = 0;
disk_mem[ 5337] = 0;
disk_mem[ 5338] = 0;
disk_mem[ 5339] = 0;
disk_mem[ 5340] = 0;
disk_mem[ 5341] = 0;
disk_mem[ 5342] = 0;
disk_mem[ 5343] = 0;
disk_mem[ 5344] = 0;
disk_mem[ 5345] = 0;
disk_mem[ 5346] = 0;
disk_mem[ 5347] = 0;
disk_mem[ 5348] = 0;
disk_mem[ 5349] = 0;
disk_mem[ 5350] = 0;
disk_mem[ 5351] = 0;
disk_mem[ 5352] = 0;
disk_mem[ 5353] = 0;
disk_mem[ 5354] = 0;
disk_mem[ 5355] = 0;
disk_mem[ 5356] = 0;
disk_mem[ 5357] = 0;
disk_mem[ 5358] = 0;
disk_mem[ 5359] = 0;
disk_mem[ 5360] = 0;
disk_mem[ 5361] = 0;
disk_mem[ 5362] = 0;
disk_mem[ 5363] = 0;
disk_mem[ 5364] = 0;
disk_mem[ 5365] = 0;
disk_mem[ 5366] = 0;
disk_mem[ 5367] = 0;
disk_mem[ 5368] = 0;
disk_mem[ 5369] = 0;
disk_mem[ 5370] = 0;
disk_mem[ 5371] = 0;
disk_mem[ 5372] = 0;
disk_mem[ 5373] = 0;
disk_mem[ 5374] = 0;
disk_mem[ 5375] = 0;
disk_mem[ 5376] = 0;
disk_mem[ 5377] = 0;
disk_mem[ 5378] = 0;
disk_mem[ 5379] = 0;
disk_mem[ 5380] = 0;
disk_mem[ 5381] = 0;
disk_mem[ 5382] = 0;
disk_mem[ 5383] = 0;
disk_mem[ 5384] = 0;
disk_mem[ 5385] = 0;
disk_mem[ 5386] = 0;
disk_mem[ 5387] = 0;
disk_mem[ 5388] = 0;
disk_mem[ 5389] = 0;
disk_mem[ 5390] = 0;
disk_mem[ 5391] = 0;
disk_mem[ 5392] = 0;
disk_mem[ 5393] = 0;
disk_mem[ 5394] = 0;
disk_mem[ 5395] = 0;
disk_mem[ 5396] = 0;
disk_mem[ 5397] = 0;
disk_mem[ 5398] = 0;
disk_mem[ 5399] = 0;
disk_mem[ 5400] = 0;
disk_mem[ 5401] = 0;
disk_mem[ 5402] = 0;
disk_mem[ 5403] = 0;
disk_mem[ 5404] = 0;
disk_mem[ 5405] = 0;
disk_mem[ 5406] = 0;
disk_mem[ 5407] = 0;
disk_mem[ 5408] = 0;
disk_mem[ 5409] = 0;
disk_mem[ 5410] = 0;
disk_mem[ 5411] = 0;
disk_mem[ 5412] = 0;
disk_mem[ 5413] = 0;
disk_mem[ 5414] = 0;
disk_mem[ 5415] = 0;
disk_mem[ 5416] = 0;
disk_mem[ 5417] = 0;
disk_mem[ 5418] = 0;
disk_mem[ 5419] = 0;
disk_mem[ 5420] = 0;
disk_mem[ 5421] = 0;
disk_mem[ 5422] = 0;
disk_mem[ 5423] = 0;
disk_mem[ 5424] = 0;
disk_mem[ 5425] = 0;
disk_mem[ 5426] = 0;
disk_mem[ 5427] = 0;
disk_mem[ 5428] = 0;
disk_mem[ 5429] = 0;
disk_mem[ 5430] = 0;
disk_mem[ 5431] = 0;
disk_mem[ 5432] = 0;
disk_mem[ 5433] = 0;
disk_mem[ 5434] = 0;
disk_mem[ 5435] = 0;
disk_mem[ 5436] = 0;
disk_mem[ 5437] = 0;
disk_mem[ 5438] = 0;
disk_mem[ 5439] = 0;
disk_mem[ 5440] = 0;
disk_mem[ 5441] = 0;
disk_mem[ 5442] = 0;
disk_mem[ 5443] = 0;
disk_mem[ 5444] = 0;
disk_mem[ 5445] = 0;
disk_mem[ 5446] = 0;
disk_mem[ 5447] = 0;
disk_mem[ 5448] = 0;
disk_mem[ 5449] = 0;
disk_mem[ 5450] = 0;
disk_mem[ 5451] = 0;
disk_mem[ 5452] = 0;
disk_mem[ 5453] = 0;
disk_mem[ 5454] = 0;
disk_mem[ 5455] = 0;
disk_mem[ 5456] = 0;
disk_mem[ 5457] = 0;
disk_mem[ 5458] = 0;
disk_mem[ 5459] = 0;
disk_mem[ 5460] = 0;
disk_mem[ 5461] = 0;
disk_mem[ 5462] = 0;
disk_mem[ 5463] = 0;
disk_mem[ 5464] = 0;
disk_mem[ 5465] = 0;
disk_mem[ 5466] = 0;
disk_mem[ 5467] = 0;
disk_mem[ 5468] = 0;
disk_mem[ 5469] = 0;
disk_mem[ 5470] = 0;
disk_mem[ 5471] = 0;
disk_mem[ 5472] = 0;
disk_mem[ 5473] = 0;
disk_mem[ 5474] = 0;
disk_mem[ 5475] = 0;
disk_mem[ 5476] = 0;
disk_mem[ 5477] = 0;
disk_mem[ 5478] = 0;
disk_mem[ 5479] = 0;
disk_mem[ 5480] = 0;
disk_mem[ 5481] = 0;
disk_mem[ 5482] = 0;
disk_mem[ 5483] = 0;
disk_mem[ 5484] = 0;
disk_mem[ 5485] = 0;
disk_mem[ 5486] = 0;
disk_mem[ 5487] = 0;
disk_mem[ 5488] = 0;
disk_mem[ 5489] = 0;
disk_mem[ 5490] = 0;
disk_mem[ 5491] = 0;
disk_mem[ 5492] = 0;
disk_mem[ 5493] = 0;
disk_mem[ 5494] = 0;
disk_mem[ 5495] = 0;
disk_mem[ 5496] = 0;
disk_mem[ 5497] = 0;
disk_mem[ 5498] = 0;
disk_mem[ 5499] = 0;
disk_mem[ 5500] = 0;
disk_mem[ 5501] = 0;
disk_mem[ 5502] = 0;
disk_mem[ 5503] = 0;
disk_mem[ 5504] = 0;
disk_mem[ 5505] = 0;
disk_mem[ 5506] = 0;
disk_mem[ 5507] = 0;
disk_mem[ 5508] = 0;
disk_mem[ 5509] = 0;
disk_mem[ 5510] = 0;
disk_mem[ 5511] = 0;
disk_mem[ 5512] = 0;
disk_mem[ 5513] = 0;
disk_mem[ 5514] = 0;
disk_mem[ 5515] = 0;
disk_mem[ 5516] = 0;
disk_mem[ 5517] = 0;
disk_mem[ 5518] = 0;
disk_mem[ 5519] = 0;
disk_mem[ 5520] = 0;
disk_mem[ 5521] = 0;
disk_mem[ 5522] = 0;
disk_mem[ 5523] = 0;
disk_mem[ 5524] = 0;
disk_mem[ 5525] = 0;
disk_mem[ 5526] = 0;
disk_mem[ 5527] = 0;
disk_mem[ 5528] = 0;
disk_mem[ 5529] = 0;
disk_mem[ 5530] = 0;
disk_mem[ 5531] = 0;
disk_mem[ 5532] = 0;
disk_mem[ 5533] = 0;
disk_mem[ 5534] = 0;
disk_mem[ 5535] = 0;
disk_mem[ 5536] = 0;
disk_mem[ 5537] = 0;
disk_mem[ 5538] = 0;
disk_mem[ 5539] = 0;
disk_mem[ 5540] = 0;
disk_mem[ 5541] = 0;
disk_mem[ 5542] = 0;
disk_mem[ 5543] = 0;
disk_mem[ 5544] = 0;
disk_mem[ 5545] = 0;
disk_mem[ 5546] = 0;
disk_mem[ 5547] = 0;
disk_mem[ 5548] = 0;
disk_mem[ 5549] = 0;
disk_mem[ 5550] = 0;
disk_mem[ 5551] = 0;
disk_mem[ 5552] = 0;
disk_mem[ 5553] = 0;
disk_mem[ 5554] = 0;
disk_mem[ 5555] = 0;
disk_mem[ 5556] = 0;
disk_mem[ 5557] = 0;
disk_mem[ 5558] = 0;
disk_mem[ 5559] = 0;
disk_mem[ 5560] = 0;
disk_mem[ 5561] = 0;
disk_mem[ 5562] = 0;
disk_mem[ 5563] = 0;
disk_mem[ 5564] = 0;
disk_mem[ 5565] = 0;
disk_mem[ 5566] = 0;
disk_mem[ 5567] = 0;
disk_mem[ 5568] = 0;
disk_mem[ 5569] = 0;
disk_mem[ 5570] = 0;
disk_mem[ 5571] = 0;
disk_mem[ 5572] = 0;
disk_mem[ 5573] = 0;
disk_mem[ 5574] = 0;
disk_mem[ 5575] = 0;
disk_mem[ 5576] = 0;
disk_mem[ 5577] = 0;
disk_mem[ 5578] = 0;
disk_mem[ 5579] = 0;
disk_mem[ 5580] = 0;
disk_mem[ 5581] = 0;
disk_mem[ 5582] = 0;
disk_mem[ 5583] = 0;
disk_mem[ 5584] = 0;
disk_mem[ 5585] = 0;
disk_mem[ 5586] = 0;
disk_mem[ 5587] = 0;
disk_mem[ 5588] = 0;
disk_mem[ 5589] = 0;
disk_mem[ 5590] = 0;
disk_mem[ 5591] = 0;
disk_mem[ 5592] = 0;
disk_mem[ 5593] = 0;
disk_mem[ 5594] = 0;
disk_mem[ 5595] = 0;
disk_mem[ 5596] = 0;
disk_mem[ 5597] = 0;
disk_mem[ 5598] = 0;
disk_mem[ 5599] = 0;
disk_mem[ 5600] = 0;
disk_mem[ 5601] = 0;
disk_mem[ 5602] = 0;
disk_mem[ 5603] = 0;
disk_mem[ 5604] = 0;
disk_mem[ 5605] = 0;
disk_mem[ 5606] = 0;
disk_mem[ 5607] = 0;
disk_mem[ 5608] = 0;
disk_mem[ 5609] = 0;
disk_mem[ 5610] = 0;
disk_mem[ 5611] = 0;
disk_mem[ 5612] = 0;
disk_mem[ 5613] = 0;
disk_mem[ 5614] = 0;
disk_mem[ 5615] = 0;
disk_mem[ 5616] = 0;
disk_mem[ 5617] = 0;
disk_mem[ 5618] = 0;
disk_mem[ 5619] = 0;
disk_mem[ 5620] = 0;
disk_mem[ 5621] = 0;
disk_mem[ 5622] = 0;
disk_mem[ 5623] = 0;
disk_mem[ 5624] = 0;
disk_mem[ 5625] = 0;
disk_mem[ 5626] = 0;
disk_mem[ 5627] = 0;
disk_mem[ 5628] = 0;
disk_mem[ 5629] = 0;
disk_mem[ 5630] = 0;
disk_mem[ 5631] = 0;
disk_mem[ 5632] = 0;
disk_mem[ 5633] = 0;
disk_mem[ 5634] = 0;
disk_mem[ 5635] = 0;
disk_mem[ 5636] = 0;
disk_mem[ 5637] = 0;
disk_mem[ 5638] = 0;
disk_mem[ 5639] = 0;
disk_mem[ 5640] = 0;
disk_mem[ 5641] = 0;
disk_mem[ 5642] = 0;
disk_mem[ 5643] = 0;
disk_mem[ 5644] = 0;
disk_mem[ 5645] = 0;
disk_mem[ 5646] = 0;
disk_mem[ 5647] = 0;
disk_mem[ 5648] = 0;
disk_mem[ 5649] = 0;
disk_mem[ 5650] = 0;
disk_mem[ 5651] = 0;
disk_mem[ 5652] = 0;
disk_mem[ 5653] = 0;
disk_mem[ 5654] = 0;
disk_mem[ 5655] = 0;
disk_mem[ 5656] = 0;
disk_mem[ 5657] = 0;
disk_mem[ 5658] = 0;
disk_mem[ 5659] = 0;
disk_mem[ 5660] = 0;
disk_mem[ 5661] = 0;
disk_mem[ 5662] = 0;
disk_mem[ 5663] = 0;
disk_mem[ 5664] = 0;
disk_mem[ 5665] = 0;
disk_mem[ 5666] = 0;
disk_mem[ 5667] = 0;
disk_mem[ 5668] = 0;
disk_mem[ 5669] = 0;
disk_mem[ 5670] = 0;
disk_mem[ 5671] = 0;
disk_mem[ 5672] = 0;
disk_mem[ 5673] = 0;
disk_mem[ 5674] = 0;
disk_mem[ 5675] = 0;
disk_mem[ 5676] = 0;
disk_mem[ 5677] = 0;
disk_mem[ 5678] = 0;
disk_mem[ 5679] = 0;
disk_mem[ 5680] = 0;
disk_mem[ 5681] = 0;
disk_mem[ 5682] = 0;
disk_mem[ 5683] = 0;
disk_mem[ 5684] = 0;
disk_mem[ 5685] = 0;
disk_mem[ 5686] = 0;
disk_mem[ 5687] = 0;
disk_mem[ 5688] = 0;
disk_mem[ 5689] = 0;
disk_mem[ 5690] = 0;
disk_mem[ 5691] = 0;
disk_mem[ 5692] = 0;
disk_mem[ 5693] = 0;
disk_mem[ 5694] = 0;
disk_mem[ 5695] = 0;
disk_mem[ 5696] = 0;
disk_mem[ 5697] = 0;
disk_mem[ 5698] = 0;
disk_mem[ 5699] = 0;
disk_mem[ 5700] = 0;
disk_mem[ 5701] = 0;
disk_mem[ 5702] = 0;
disk_mem[ 5703] = 0;
disk_mem[ 5704] = 0;
disk_mem[ 5705] = 0;
disk_mem[ 5706] = 0;
disk_mem[ 5707] = 0;
disk_mem[ 5708] = 0;
disk_mem[ 5709] = 0;
disk_mem[ 5710] = 0;
disk_mem[ 5711] = 0;
disk_mem[ 5712] = 0;
disk_mem[ 5713] = 0;
disk_mem[ 5714] = 0;
disk_mem[ 5715] = 0;
disk_mem[ 5716] = 0;
disk_mem[ 5717] = 0;
disk_mem[ 5718] = 0;
disk_mem[ 5719] = 0;
disk_mem[ 5720] = 0;
disk_mem[ 5721] = 0;
disk_mem[ 5722] = 0;
disk_mem[ 5723] = 0;
disk_mem[ 5724] = 0;
disk_mem[ 5725] = 0;
disk_mem[ 5726] = 0;
disk_mem[ 5727] = 0;
disk_mem[ 5728] = 0;
disk_mem[ 5729] = 0;
disk_mem[ 5730] = 0;
disk_mem[ 5731] = 0;
disk_mem[ 5732] = 0;
disk_mem[ 5733] = 0;
disk_mem[ 5734] = 0;
disk_mem[ 5735] = 0;
disk_mem[ 5736] = 0;
disk_mem[ 5737] = 0;
disk_mem[ 5738] = 0;
disk_mem[ 5739] = 0;
disk_mem[ 5740] = 0;
disk_mem[ 5741] = 0;
disk_mem[ 5742] = 0;
disk_mem[ 5743] = 0;
disk_mem[ 5744] = 0;
disk_mem[ 5745] = 0;
disk_mem[ 5746] = 0;
disk_mem[ 5747] = 0;
disk_mem[ 5748] = 0;
disk_mem[ 5749] = 0;
disk_mem[ 5750] = 0;
disk_mem[ 5751] = 0;
disk_mem[ 5752] = 0;
disk_mem[ 5753] = 0;
disk_mem[ 5754] = 0;
disk_mem[ 5755] = 0;
disk_mem[ 5756] = 0;
disk_mem[ 5757] = 0;
disk_mem[ 5758] = 0;
disk_mem[ 5759] = 0;
disk_mem[ 5760] = 0;
disk_mem[ 5761] = 0;
disk_mem[ 5762] = 0;
disk_mem[ 5763] = 0;
disk_mem[ 5764] = 0;
disk_mem[ 5765] = 0;
disk_mem[ 5766] = 0;
disk_mem[ 5767] = 0;
disk_mem[ 5768] = 0;
disk_mem[ 5769] = 0;
disk_mem[ 5770] = 0;
disk_mem[ 5771] = 0;
disk_mem[ 5772] = 0;
disk_mem[ 5773] = 0;
disk_mem[ 5774] = 0;
disk_mem[ 5775] = 0;
disk_mem[ 5776] = 0;
disk_mem[ 5777] = 0;
disk_mem[ 5778] = 0;
disk_mem[ 5779] = 0;
disk_mem[ 5780] = 0;
disk_mem[ 5781] = 0;
disk_mem[ 5782] = 0;
disk_mem[ 5783] = 0;
disk_mem[ 5784] = 0;
disk_mem[ 5785] = 0;
disk_mem[ 5786] = 0;
disk_mem[ 5787] = 0;
disk_mem[ 5788] = 0;
disk_mem[ 5789] = 0;
disk_mem[ 5790] = 0;
disk_mem[ 5791] = 0;
disk_mem[ 5792] = 0;
disk_mem[ 5793] = 0;
disk_mem[ 5794] = 0;
disk_mem[ 5795] = 0;
disk_mem[ 5796] = 0;
disk_mem[ 5797] = 0;
disk_mem[ 5798] = 0;
disk_mem[ 5799] = 0;
disk_mem[ 5800] = 0;
disk_mem[ 5801] = 0;
disk_mem[ 5802] = 0;
disk_mem[ 5803] = 0;
disk_mem[ 5804] = 0;
disk_mem[ 5805] = 0;
disk_mem[ 5806] = 0;
disk_mem[ 5807] = 0;
disk_mem[ 5808] = 0;
disk_mem[ 5809] = 0;
disk_mem[ 5810] = 0;
disk_mem[ 5811] = 0;
disk_mem[ 5812] = 0;
disk_mem[ 5813] = 0;
disk_mem[ 5814] = 0;
disk_mem[ 5815] = 0;
disk_mem[ 5816] = 0;
disk_mem[ 5817] = 0;
disk_mem[ 5818] = 0;
disk_mem[ 5819] = 0;
disk_mem[ 5820] = 0;
disk_mem[ 5821] = 0;
disk_mem[ 5822] = 0;
disk_mem[ 5823] = 0;
disk_mem[ 5824] = 0;
disk_mem[ 5825] = 0;
disk_mem[ 5826] = 0;
disk_mem[ 5827] = 0;
disk_mem[ 5828] = 0;
disk_mem[ 5829] = 0;
disk_mem[ 5830] = 0;
disk_mem[ 5831] = 0;
disk_mem[ 5832] = 0;
disk_mem[ 5833] = 0;
disk_mem[ 5834] = 0;
disk_mem[ 5835] = 0;
disk_mem[ 5836] = 0;
disk_mem[ 5837] = 0;
disk_mem[ 5838] = 0;
disk_mem[ 5839] = 0;
disk_mem[ 5840] = 0;
disk_mem[ 5841] = 0;
disk_mem[ 5842] = 0;
disk_mem[ 5843] = 0;
disk_mem[ 5844] = 0;
disk_mem[ 5845] = 0;
disk_mem[ 5846] = 0;
disk_mem[ 5847] = 0;
disk_mem[ 5848] = 0;
disk_mem[ 5849] = 0;
disk_mem[ 5850] = 0;
disk_mem[ 5851] = 0;
disk_mem[ 5852] = 0;
disk_mem[ 5853] = 0;
disk_mem[ 5854] = 0;
disk_mem[ 5855] = 0;
disk_mem[ 5856] = 0;
disk_mem[ 5857] = 0;
disk_mem[ 5858] = 0;
disk_mem[ 5859] = 0;
disk_mem[ 5860] = 0;
disk_mem[ 5861] = 0;
disk_mem[ 5862] = 0;
disk_mem[ 5863] = 0;
disk_mem[ 5864] = 0;
disk_mem[ 5865] = 0;
disk_mem[ 5866] = 0;
disk_mem[ 5867] = 0;
disk_mem[ 5868] = 0;
disk_mem[ 5869] = 0;
disk_mem[ 5870] = 0;
disk_mem[ 5871] = 0;
disk_mem[ 5872] = 0;
disk_mem[ 5873] = 0;
disk_mem[ 5874] = 0;
disk_mem[ 5875] = 0;
disk_mem[ 5876] = 0;
disk_mem[ 5877] = 0;
disk_mem[ 5878] = 0;
disk_mem[ 5879] = 0;
disk_mem[ 5880] = 0;
disk_mem[ 5881] = 0;
disk_mem[ 5882] = 0;
disk_mem[ 5883] = 0;
disk_mem[ 5884] = 0;
disk_mem[ 5885] = 0;
disk_mem[ 5886] = 0;
disk_mem[ 5887] = 0;
disk_mem[ 5888] = 0;
disk_mem[ 5889] = 0;
disk_mem[ 5890] = 0;
disk_mem[ 5891] = 0;
disk_mem[ 5892] = 0;
disk_mem[ 5893] = 0;
disk_mem[ 5894] = 0;
disk_mem[ 5895] = 0;
disk_mem[ 5896] = 0;
disk_mem[ 5897] = 0;
disk_mem[ 5898] = 0;
disk_mem[ 5899] = 0;
disk_mem[ 5900] = 0;
disk_mem[ 5901] = 0;
disk_mem[ 5902] = 0;
disk_mem[ 5903] = 0;
disk_mem[ 5904] = 0;
disk_mem[ 5905] = 0;
disk_mem[ 5906] = 0;
disk_mem[ 5907] = 0;
disk_mem[ 5908] = 0;
disk_mem[ 5909] = 0;
disk_mem[ 5910] = 0;
disk_mem[ 5911] = 0;
disk_mem[ 5912] = 0;
disk_mem[ 5913] = 0;
disk_mem[ 5914] = 0;
disk_mem[ 5915] = 0;
disk_mem[ 5916] = 0;
disk_mem[ 5917] = 0;
disk_mem[ 5918] = 0;
disk_mem[ 5919] = 0;
disk_mem[ 5920] = 0;
disk_mem[ 5921] = 0;
disk_mem[ 5922] = 0;
disk_mem[ 5923] = 0;
disk_mem[ 5924] = 0;
disk_mem[ 5925] = 0;
disk_mem[ 5926] = 0;
disk_mem[ 5927] = 0;
disk_mem[ 5928] = 0;
disk_mem[ 5929] = 0;
disk_mem[ 5930] = 0;
disk_mem[ 5931] = 0;
disk_mem[ 5932] = 0;
disk_mem[ 5933] = 0;
disk_mem[ 5934] = 0;
disk_mem[ 5935] = 0;
disk_mem[ 5936] = 0;
disk_mem[ 5937] = 0;
disk_mem[ 5938] = 0;
disk_mem[ 5939] = 0;
disk_mem[ 5940] = 0;
disk_mem[ 5941] = 0;
disk_mem[ 5942] = 0;
disk_mem[ 5943] = 0;
disk_mem[ 5944] = 0;
disk_mem[ 5945] = 0;
disk_mem[ 5946] = 0;
disk_mem[ 5947] = 0;
disk_mem[ 5948] = 0;
disk_mem[ 5949] = 0;
disk_mem[ 5950] = 0;
disk_mem[ 5951] = 0;
disk_mem[ 5952] = 0;
disk_mem[ 5953] = 0;
disk_mem[ 5954] = 0;
disk_mem[ 5955] = 0;
disk_mem[ 5956] = 0;
disk_mem[ 5957] = 0;
disk_mem[ 5958] = 0;
disk_mem[ 5959] = 0;
disk_mem[ 5960] = 0;
disk_mem[ 5961] = 0;
disk_mem[ 5962] = 0;
disk_mem[ 5963] = 0;
disk_mem[ 5964] = 0;
disk_mem[ 5965] = 0;
disk_mem[ 5966] = 0;
disk_mem[ 5967] = 0;
disk_mem[ 5968] = 0;
disk_mem[ 5969] = 0;
disk_mem[ 5970] = 0;
disk_mem[ 5971] = 0;
disk_mem[ 5972] = 0;
disk_mem[ 5973] = 0;
disk_mem[ 5974] = 0;
disk_mem[ 5975] = 0;
disk_mem[ 5976] = 0;
disk_mem[ 5977] = 0;
disk_mem[ 5978] = 0;
disk_mem[ 5979] = 0;
disk_mem[ 5980] = 0;
disk_mem[ 5981] = 0;
disk_mem[ 5982] = 0;
disk_mem[ 5983] = 0;
disk_mem[ 5984] = 0;
disk_mem[ 5985] = 0;
disk_mem[ 5986] = 0;
disk_mem[ 5987] = 0;
disk_mem[ 5988] = 0;
disk_mem[ 5989] = 0;
disk_mem[ 5990] = 0;
disk_mem[ 5991] = 0;
disk_mem[ 5992] = 0;
disk_mem[ 5993] = 0;
disk_mem[ 5994] = 0;
disk_mem[ 5995] = 0;
disk_mem[ 5996] = 0;
disk_mem[ 5997] = 0;
disk_mem[ 5998] = 0;
disk_mem[ 5999] = 0;
disk_mem[ 6000] = 0;
disk_mem[ 6001] = 0;
disk_mem[ 6002] = 0;
disk_mem[ 6003] = 0;
disk_mem[ 6004] = 0;
disk_mem[ 6005] = 0;
disk_mem[ 6006] = 0;
disk_mem[ 6007] = 0;
disk_mem[ 6008] = 0;
disk_mem[ 6009] = 0;
disk_mem[ 6010] = 0;
disk_mem[ 6011] = 0;
disk_mem[ 6012] = 0;
disk_mem[ 6013] = 0;
disk_mem[ 6014] = 0;
disk_mem[ 6015] = 0;
disk_mem[ 6016] = 0;
disk_mem[ 6017] = 0;
disk_mem[ 6018] = 0;
disk_mem[ 6019] = 0;
disk_mem[ 6020] = 0;
disk_mem[ 6021] = 0;
disk_mem[ 6022] = 0;
disk_mem[ 6023] = 0;
disk_mem[ 6024] = 0;
disk_mem[ 6025] = 0;
disk_mem[ 6026] = 0;
disk_mem[ 6027] = 0;
disk_mem[ 6028] = 0;
disk_mem[ 6029] = 0;
disk_mem[ 6030] = 0;
disk_mem[ 6031] = 0;
disk_mem[ 6032] = 0;
disk_mem[ 6033] = 0;
disk_mem[ 6034] = 0;
disk_mem[ 6035] = 0;
disk_mem[ 6036] = 0;
disk_mem[ 6037] = 0;
disk_mem[ 6038] = 0;
disk_mem[ 6039] = 0;
disk_mem[ 6040] = 0;
disk_mem[ 6041] = 0;
disk_mem[ 6042] = 0;
disk_mem[ 6043] = 0;
disk_mem[ 6044] = 0;
disk_mem[ 6045] = 0;
disk_mem[ 6046] = 0;
disk_mem[ 6047] = 0;
disk_mem[ 6048] = 0;
disk_mem[ 6049] = 0;
disk_mem[ 6050] = 0;
disk_mem[ 6051] = 0;
disk_mem[ 6052] = 0;
disk_mem[ 6053] = 0;
disk_mem[ 6054] = 0;
disk_mem[ 6055] = 0;
disk_mem[ 6056] = 0;
disk_mem[ 6057] = 0;
disk_mem[ 6058] = 0;
disk_mem[ 6059] = 0;
disk_mem[ 6060] = 0;
disk_mem[ 6061] = 0;
disk_mem[ 6062] = 0;
disk_mem[ 6063] = 0;
disk_mem[ 6064] = 0;
disk_mem[ 6065] = 0;
disk_mem[ 6066] = 0;
disk_mem[ 6067] = 0;
disk_mem[ 6068] = 0;
disk_mem[ 6069] = 0;
disk_mem[ 6070] = 0;
disk_mem[ 6071] = 0;
disk_mem[ 6072] = 0;
disk_mem[ 6073] = 0;
disk_mem[ 6074] = 0;
disk_mem[ 6075] = 0;
disk_mem[ 6076] = 0;
disk_mem[ 6077] = 0;
disk_mem[ 6078] = 0;
disk_mem[ 6079] = 0;
disk_mem[ 6080] = 0;
disk_mem[ 6081] = 0;
disk_mem[ 6082] = 0;
disk_mem[ 6083] = 0;
disk_mem[ 6084] = 0;
disk_mem[ 6085] = 0;
disk_mem[ 6086] = 0;
disk_mem[ 6087] = 0;
disk_mem[ 6088] = 0;
disk_mem[ 6089] = 0;
disk_mem[ 6090] = 0;
disk_mem[ 6091] = 0;
disk_mem[ 6092] = 0;
disk_mem[ 6093] = 0;
disk_mem[ 6094] = 0;
disk_mem[ 6095] = 0;
disk_mem[ 6096] = 0;
disk_mem[ 6097] = 0;
disk_mem[ 6098] = 0;
disk_mem[ 6099] = 0;
disk_mem[ 6100] = 0;
disk_mem[ 6101] = 0;
disk_mem[ 6102] = 0;
disk_mem[ 6103] = 0;
disk_mem[ 6104] = 0;
disk_mem[ 6105] = 0;
disk_mem[ 6106] = 0;
disk_mem[ 6107] = 0;
disk_mem[ 6108] = 0;
disk_mem[ 6109] = 0;
disk_mem[ 6110] = 0;
disk_mem[ 6111] = 0;
disk_mem[ 6112] = 0;
disk_mem[ 6113] = 0;
disk_mem[ 6114] = 0;
disk_mem[ 6115] = 0;
disk_mem[ 6116] = 0;
disk_mem[ 6117] = 0;
disk_mem[ 6118] = 0;
disk_mem[ 6119] = 0;
disk_mem[ 6120] = 0;
disk_mem[ 6121] = 0;
disk_mem[ 6122] = 0;
disk_mem[ 6123] = 0;
disk_mem[ 6124] = 0;
disk_mem[ 6125] = 0;
disk_mem[ 6126] = 0;
disk_mem[ 6127] = 0;
disk_mem[ 6128] = 0;
disk_mem[ 6129] = 0;
disk_mem[ 6130] = 0;
disk_mem[ 6131] = 0;
disk_mem[ 6132] = 0;
disk_mem[ 6133] = 0;
disk_mem[ 6134] = 0;
disk_mem[ 6135] = 0;
disk_mem[ 6136] = 0;
disk_mem[ 6137] = 0;
disk_mem[ 6138] = 0;
disk_mem[ 6139] = 0;
disk_mem[ 6140] = 0;
disk_mem[ 6141] = 0;
disk_mem[ 6142] = 0;
disk_mem[ 6143] = 0;
disk_mem[ 6144] = 0;
disk_mem[ 6145] = 0;
disk_mem[ 6146] = 0;
disk_mem[ 6147] = 0;
disk_mem[ 6148] = 0;
disk_mem[ 6149] = 0;
disk_mem[ 6150] = 0;
disk_mem[ 6151] = 0;
disk_mem[ 6152] = 0;
disk_mem[ 6153] = 0;
disk_mem[ 6154] = 0;
disk_mem[ 6155] = 0;
disk_mem[ 6156] = 0;
disk_mem[ 6157] = 0;
disk_mem[ 6158] = 0;
disk_mem[ 6159] = 0;
disk_mem[ 6160] = 0;
disk_mem[ 6161] = 0;
disk_mem[ 6162] = 0;
disk_mem[ 6163] = 0;
disk_mem[ 6164] = 0;
disk_mem[ 6165] = 0;
disk_mem[ 6166] = 0;
disk_mem[ 6167] = 0;
disk_mem[ 6168] = 0;
disk_mem[ 6169] = 0;
disk_mem[ 6170] = 0;
disk_mem[ 6171] = 0;
disk_mem[ 6172] = 0;
disk_mem[ 6173] = 0;
disk_mem[ 6174] = 0;
disk_mem[ 6175] = 0;
disk_mem[ 6176] = 0;
disk_mem[ 6177] = 0;
disk_mem[ 6178] = 0;
disk_mem[ 6179] = 0;
disk_mem[ 6180] = 0;
disk_mem[ 6181] = 0;
disk_mem[ 6182] = 0;
disk_mem[ 6183] = 0;
disk_mem[ 6184] = 0;
disk_mem[ 6185] = 0;
disk_mem[ 6186] = 0;
disk_mem[ 6187] = 0;
disk_mem[ 6188] = 0;
disk_mem[ 6189] = 0;
disk_mem[ 6190] = 0;
disk_mem[ 6191] = 0;
disk_mem[ 6192] = 0;
disk_mem[ 6193] = 0;
disk_mem[ 6194] = 0;
disk_mem[ 6195] = 0;
disk_mem[ 6196] = 0;
disk_mem[ 6197] = 0;
disk_mem[ 6198] = 0;
disk_mem[ 6199] = 0;
disk_mem[ 6200] = 0;
disk_mem[ 6201] = 0;
disk_mem[ 6202] = 0;
disk_mem[ 6203] = 0;
disk_mem[ 6204] = 0;
disk_mem[ 6205] = 0;
disk_mem[ 6206] = 0;
disk_mem[ 6207] = 0;
disk_mem[ 6208] = 0;
disk_mem[ 6209] = 0;
disk_mem[ 6210] = 0;
disk_mem[ 6211] = 0;
disk_mem[ 6212] = 0;
disk_mem[ 6213] = 0;
disk_mem[ 6214] = 0;
disk_mem[ 6215] = 0;
disk_mem[ 6216] = 0;
disk_mem[ 6217] = 0;
disk_mem[ 6218] = 0;
disk_mem[ 6219] = 0;
disk_mem[ 6220] = 0;
disk_mem[ 6221] = 0;
disk_mem[ 6222] = 0;
disk_mem[ 6223] = 0;
disk_mem[ 6224] = 0;
disk_mem[ 6225] = 0;
disk_mem[ 6226] = 0;
disk_mem[ 6227] = 0;
disk_mem[ 6228] = 0;
disk_mem[ 6229] = 0;
disk_mem[ 6230] = 0;
disk_mem[ 6231] = 0;
disk_mem[ 6232] = 0;
disk_mem[ 6233] = 0;
disk_mem[ 6234] = 0;
disk_mem[ 6235] = 0;
disk_mem[ 6236] = 0;
disk_mem[ 6237] = 0;
disk_mem[ 6238] = 0;
disk_mem[ 6239] = 0;
disk_mem[ 6240] = 0;
disk_mem[ 6241] = 0;
disk_mem[ 6242] = 0;
disk_mem[ 6243] = 0;
disk_mem[ 6244] = 0;
disk_mem[ 6245] = 0;
disk_mem[ 6246] = 0;
disk_mem[ 6247] = 0;
disk_mem[ 6248] = 0;
disk_mem[ 6249] = 0;
disk_mem[ 6250] = 0;
disk_mem[ 6251] = 0;
disk_mem[ 6252] = 0;
disk_mem[ 6253] = 0;
disk_mem[ 6254] = 0;
disk_mem[ 6255] = 0;
disk_mem[ 6256] = 0;
disk_mem[ 6257] = 0;
disk_mem[ 6258] = 0;
disk_mem[ 6259] = 0;
disk_mem[ 6260] = 0;
disk_mem[ 6261] = 0;
disk_mem[ 6262] = 0;
disk_mem[ 6263] = 0;
disk_mem[ 6264] = 0;
disk_mem[ 6265] = 0;
disk_mem[ 6266] = 0;
disk_mem[ 6267] = 0;
disk_mem[ 6268] = 0;
disk_mem[ 6269] = 0;
disk_mem[ 6270] = 0;
disk_mem[ 6271] = 0;
disk_mem[ 6272] = 0;
disk_mem[ 6273] = 0;
disk_mem[ 6274] = 0;
disk_mem[ 6275] = 0;
disk_mem[ 6276] = 0;
disk_mem[ 6277] = 0;
disk_mem[ 6278] = 0;
disk_mem[ 6279] = 0;
disk_mem[ 6280] = 0;
disk_mem[ 6281] = 0;
disk_mem[ 6282] = 0;
disk_mem[ 6283] = 0;
disk_mem[ 6284] = 0;
disk_mem[ 6285] = 0;
disk_mem[ 6286] = 0;
disk_mem[ 6287] = 0;
disk_mem[ 6288] = 0;
disk_mem[ 6289] = 0;
disk_mem[ 6290] = 0;
disk_mem[ 6291] = 0;
disk_mem[ 6292] = 0;
disk_mem[ 6293] = 0;
disk_mem[ 6294] = 0;
disk_mem[ 6295] = 0;
disk_mem[ 6296] = 0;
disk_mem[ 6297] = 0;
disk_mem[ 6298] = 0;
disk_mem[ 6299] = 0;
disk_mem[ 6300] = 0;
disk_mem[ 6301] = 0;
disk_mem[ 6302] = 0;
disk_mem[ 6303] = 0;
disk_mem[ 6304] = 0;
disk_mem[ 6305] = 0;
disk_mem[ 6306] = 0;
disk_mem[ 6307] = 0;
disk_mem[ 6308] = 0;
disk_mem[ 6309] = 0;
disk_mem[ 6310] = 0;
disk_mem[ 6311] = 0;
disk_mem[ 6312] = 0;
disk_mem[ 6313] = 0;
disk_mem[ 6314] = 0;
disk_mem[ 6315] = 0;
disk_mem[ 6316] = 0;
disk_mem[ 6317] = 0;
disk_mem[ 6318] = 0;
disk_mem[ 6319] = 0;
disk_mem[ 6320] = 0;
disk_mem[ 6321] = 0;
disk_mem[ 6322] = 0;
disk_mem[ 6323] = 0;
disk_mem[ 6324] = 0;
disk_mem[ 6325] = 0;
disk_mem[ 6326] = 0;
disk_mem[ 6327] = 0;
disk_mem[ 6328] = 0;
disk_mem[ 6329] = 0;
disk_mem[ 6330] = 0;
disk_mem[ 6331] = 0;
disk_mem[ 6332] = 0;
disk_mem[ 6333] = 0;
disk_mem[ 6334] = 0;
disk_mem[ 6335] = 0;
disk_mem[ 6336] = 0;
disk_mem[ 6337] = 0;
disk_mem[ 6338] = 0;
disk_mem[ 6339] = 0;
disk_mem[ 6340] = 0;
disk_mem[ 6341] = 0;
disk_mem[ 6342] = 0;
disk_mem[ 6343] = 0;
disk_mem[ 6344] = 0;
disk_mem[ 6345] = 0;
disk_mem[ 6346] = 0;
disk_mem[ 6347] = 0;
disk_mem[ 6348] = 0;
disk_mem[ 6349] = 0;
disk_mem[ 6350] = 0;
disk_mem[ 6351] = 0;
disk_mem[ 6352] = 0;
disk_mem[ 6353] = 0;
disk_mem[ 6354] = 0;
disk_mem[ 6355] = 0;
disk_mem[ 6356] = 0;
disk_mem[ 6357] = 0;
disk_mem[ 6358] = 0;
disk_mem[ 6359] = 0;
disk_mem[ 6360] = 0;
disk_mem[ 6361] = 0;
disk_mem[ 6362] = 0;
disk_mem[ 6363] = 0;
disk_mem[ 6364] = 0;
disk_mem[ 6365] = 0;
disk_mem[ 6366] = 0;
disk_mem[ 6367] = 0;
disk_mem[ 6368] = 0;
disk_mem[ 6369] = 0;
disk_mem[ 6370] = 0;
disk_mem[ 6371] = 0;
disk_mem[ 6372] = 0;
disk_mem[ 6373] = 0;
disk_mem[ 6374] = 0;
disk_mem[ 6375] = 0;
disk_mem[ 6376] = 0;
disk_mem[ 6377] = 0;
disk_mem[ 6378] = 0;
disk_mem[ 6379] = 0;
disk_mem[ 6380] = 0;
disk_mem[ 6381] = 0;
disk_mem[ 6382] = 0;
disk_mem[ 6383] = 0;
disk_mem[ 6384] = 0;
disk_mem[ 6385] = 0;
disk_mem[ 6386] = 0;
disk_mem[ 6387] = 0;
disk_mem[ 6388] = 0;
disk_mem[ 6389] = 0;
disk_mem[ 6390] = 0;
disk_mem[ 6391] = 0;
disk_mem[ 6392] = 0;
disk_mem[ 6393] = 0;
disk_mem[ 6394] = 0;
disk_mem[ 6395] = 0;
disk_mem[ 6396] = 0;
disk_mem[ 6397] = 0;
disk_mem[ 6398] = 0;
disk_mem[ 6399] = 0;
disk_mem[ 6400] = 0;
disk_mem[ 6401] = 0;
disk_mem[ 6402] = 0;
disk_mem[ 6403] = 0;
disk_mem[ 6404] = 0;
disk_mem[ 6405] = 0;
disk_mem[ 6406] = 0;
disk_mem[ 6407] = 0;
disk_mem[ 6408] = 0;
disk_mem[ 6409] = 0;
disk_mem[ 6410] = 0;
disk_mem[ 6411] = 0;
disk_mem[ 6412] = 0;
disk_mem[ 6413] = 0;
disk_mem[ 6414] = 0;
disk_mem[ 6415] = 0;
disk_mem[ 6416] = 0;
disk_mem[ 6417] = 0;
disk_mem[ 6418] = 0;
disk_mem[ 6419] = 0;
disk_mem[ 6420] = 0;
disk_mem[ 6421] = 0;
disk_mem[ 6422] = 0;
disk_mem[ 6423] = 0;
disk_mem[ 6424] = 0;
disk_mem[ 6425] = 0;
disk_mem[ 6426] = 0;
disk_mem[ 6427] = 0;
disk_mem[ 6428] = 0;
disk_mem[ 6429] = 0;
disk_mem[ 6430] = 0;
disk_mem[ 6431] = 0;
disk_mem[ 6432] = 0;
disk_mem[ 6433] = 0;
disk_mem[ 6434] = 0;
disk_mem[ 6435] = 0;
disk_mem[ 6436] = 0;
disk_mem[ 6437] = 0;
disk_mem[ 6438] = 0;
disk_mem[ 6439] = 0;
disk_mem[ 6440] = 0;
disk_mem[ 6441] = 0;
disk_mem[ 6442] = 0;
disk_mem[ 6443] = 0;
disk_mem[ 6444] = 0;
disk_mem[ 6445] = 0;
disk_mem[ 6446] = 0;
disk_mem[ 6447] = 0;
disk_mem[ 6448] = 0;
disk_mem[ 6449] = 0;
disk_mem[ 6450] = 0;
disk_mem[ 6451] = 0;
disk_mem[ 6452] = 0;
disk_mem[ 6453] = 0;
disk_mem[ 6454] = 0;
disk_mem[ 6455] = 0;
disk_mem[ 6456] = 0;
disk_mem[ 6457] = 0;
disk_mem[ 6458] = 0;
disk_mem[ 6459] = 0;
disk_mem[ 6460] = 0;
disk_mem[ 6461] = 0;
disk_mem[ 6462] = 0;
disk_mem[ 6463] = 0;
disk_mem[ 6464] = 0;
disk_mem[ 6465] = 0;
disk_mem[ 6466] = 0;
disk_mem[ 6467] = 0;
disk_mem[ 6468] = 0;
disk_mem[ 6469] = 0;
disk_mem[ 6470] = 0;
disk_mem[ 6471] = 0;
disk_mem[ 6472] = 0;
disk_mem[ 6473] = 0;
disk_mem[ 6474] = 0;
disk_mem[ 6475] = 0;
disk_mem[ 6476] = 0;
disk_mem[ 6477] = 0;
disk_mem[ 6478] = 0;
disk_mem[ 6479] = 0;
disk_mem[ 6480] = 0;
disk_mem[ 6481] = 0;
disk_mem[ 6482] = 0;
disk_mem[ 6483] = 0;
disk_mem[ 6484] = 0;
disk_mem[ 6485] = 0;
disk_mem[ 6486] = 0;
disk_mem[ 6487] = 0;
disk_mem[ 6488] = 0;
disk_mem[ 6489] = 0;
disk_mem[ 6490] = 0;
disk_mem[ 6491] = 0;
disk_mem[ 6492] = 0;
disk_mem[ 6493] = 0;
disk_mem[ 6494] = 0;
disk_mem[ 6495] = 0;
disk_mem[ 6496] = 0;
disk_mem[ 6497] = 0;
disk_mem[ 6498] = 0;
disk_mem[ 6499] = 0;
disk_mem[ 6500] = 0;
disk_mem[ 6501] = 0;
disk_mem[ 6502] = 0;
disk_mem[ 6503] = 0;
disk_mem[ 6504] = 0;
disk_mem[ 6505] = 0;
disk_mem[ 6506] = 0;
disk_mem[ 6507] = 0;
disk_mem[ 6508] = 0;
disk_mem[ 6509] = 0;
disk_mem[ 6510] = 0;
disk_mem[ 6511] = 0;
disk_mem[ 6512] = 0;
disk_mem[ 6513] = 0;
disk_mem[ 6514] = 0;
disk_mem[ 6515] = 0;
disk_mem[ 6516] = 0;
disk_mem[ 6517] = 0;
disk_mem[ 6518] = 0;
disk_mem[ 6519] = 0;
disk_mem[ 6520] = 0;
disk_mem[ 6521] = 0;
disk_mem[ 6522] = 0;
disk_mem[ 6523] = 0;
disk_mem[ 6524] = 0;
disk_mem[ 6525] = 0;
disk_mem[ 6526] = 0;
disk_mem[ 6527] = 0;
disk_mem[ 6528] = 0;
disk_mem[ 6529] = 0;
disk_mem[ 6530] = 0;
disk_mem[ 6531] = 0;
disk_mem[ 6532] = 0;
disk_mem[ 6533] = 0;
disk_mem[ 6534] = 0;
disk_mem[ 6535] = 0;
disk_mem[ 6536] = 0;
disk_mem[ 6537] = 0;
disk_mem[ 6538] = 0;
disk_mem[ 6539] = 0;
disk_mem[ 6540] = 0;
disk_mem[ 6541] = 0;
disk_mem[ 6542] = 0;
disk_mem[ 6543] = 0;
disk_mem[ 6544] = 0;
disk_mem[ 6545] = 0;
disk_mem[ 6546] = 0;
disk_mem[ 6547] = 0;
disk_mem[ 6548] = 0;
disk_mem[ 6549] = 0;
disk_mem[ 6550] = 0;
disk_mem[ 6551] = 0;
disk_mem[ 6552] = 0;
disk_mem[ 6553] = 0;
disk_mem[ 6554] = 0;
disk_mem[ 6555] = 0;
disk_mem[ 6556] = 0;
disk_mem[ 6557] = 0;
disk_mem[ 6558] = 0;
disk_mem[ 6559] = 0;
disk_mem[ 6560] = 0;
disk_mem[ 6561] = 0;
disk_mem[ 6562] = 0;
disk_mem[ 6563] = 0;
disk_mem[ 6564] = 0;
disk_mem[ 6565] = 0;
disk_mem[ 6566] = 0;
disk_mem[ 6567] = 0;
disk_mem[ 6568] = 0;
disk_mem[ 6569] = 0;
disk_mem[ 6570] = 0;
disk_mem[ 6571] = 0;
disk_mem[ 6572] = 0;
disk_mem[ 6573] = 0;
disk_mem[ 6574] = 0;
disk_mem[ 6575] = 0;
disk_mem[ 6576] = 0;
disk_mem[ 6577] = 0;
disk_mem[ 6578] = 0;
disk_mem[ 6579] = 0;
disk_mem[ 6580] = 0;
disk_mem[ 6581] = 0;
disk_mem[ 6582] = 0;
disk_mem[ 6583] = 0;
disk_mem[ 6584] = 0;
disk_mem[ 6585] = 0;
disk_mem[ 6586] = 0;
disk_mem[ 6587] = 0;
disk_mem[ 6588] = 0;
disk_mem[ 6589] = 0;
disk_mem[ 6590] = 0;
disk_mem[ 6591] = 0;
disk_mem[ 6592] = 0;
disk_mem[ 6593] = 0;
disk_mem[ 6594] = 0;
disk_mem[ 6595] = 0;
disk_mem[ 6596] = 0;
disk_mem[ 6597] = 0;
disk_mem[ 6598] = 0;
disk_mem[ 6599] = 0;
disk_mem[ 6600] = 0;
disk_mem[ 6601] = 0;
disk_mem[ 6602] = 0;
disk_mem[ 6603] = 0;
disk_mem[ 6604] = 0;
disk_mem[ 6605] = 0;
disk_mem[ 6606] = 0;
disk_mem[ 6607] = 0;
disk_mem[ 6608] = 0;
disk_mem[ 6609] = 0;
disk_mem[ 6610] = 0;
disk_mem[ 6611] = 0;
disk_mem[ 6612] = 0;
disk_mem[ 6613] = 0;
disk_mem[ 6614] = 0;
disk_mem[ 6615] = 0;
disk_mem[ 6616] = 0;
disk_mem[ 6617] = 0;
disk_mem[ 6618] = 0;
disk_mem[ 6619] = 0;
disk_mem[ 6620] = 0;
disk_mem[ 6621] = 0;
disk_mem[ 6622] = 0;
disk_mem[ 6623] = 0;
disk_mem[ 6624] = 0;
disk_mem[ 6625] = 0;
disk_mem[ 6626] = 0;
disk_mem[ 6627] = 0;
disk_mem[ 6628] = 0;
disk_mem[ 6629] = 0;
disk_mem[ 6630] = 0;
disk_mem[ 6631] = 0;
disk_mem[ 6632] = 0;
disk_mem[ 6633] = 0;
disk_mem[ 6634] = 0;
disk_mem[ 6635] = 0;
disk_mem[ 6636] = 0;
disk_mem[ 6637] = 0;
disk_mem[ 6638] = 0;
disk_mem[ 6639] = 0;
disk_mem[ 6640] = 0;
disk_mem[ 6641] = 0;
disk_mem[ 6642] = 0;
disk_mem[ 6643] = 0;
disk_mem[ 6644] = 0;
disk_mem[ 6645] = 0;
disk_mem[ 6646] = 0;
disk_mem[ 6647] = 0;
disk_mem[ 6648] = 0;
disk_mem[ 6649] = 0;
disk_mem[ 6650] = 0;
disk_mem[ 6651] = 0;
disk_mem[ 6652] = 0;
disk_mem[ 6653] = 0;
disk_mem[ 6654] = 0;
disk_mem[ 6655] = 0;
disk_mem[ 6656] = 0;
disk_mem[ 6657] = 0;
disk_mem[ 6658] = 0;
disk_mem[ 6659] = 0;
disk_mem[ 6660] = 0;
disk_mem[ 6661] = 0;
disk_mem[ 6662] = 0;
disk_mem[ 6663] = 0;
disk_mem[ 6664] = 0;
disk_mem[ 6665] = 0;
disk_mem[ 6666] = 0;
disk_mem[ 6667] = 0;
disk_mem[ 6668] = 0;
disk_mem[ 6669] = 0;
disk_mem[ 6670] = 0;
disk_mem[ 6671] = 0;
disk_mem[ 6672] = 0;
disk_mem[ 6673] = 0;
disk_mem[ 6674] = 0;
disk_mem[ 6675] = 0;
disk_mem[ 6676] = 0;
disk_mem[ 6677] = 0;
disk_mem[ 6678] = 0;
disk_mem[ 6679] = 0;
disk_mem[ 6680] = 0;
disk_mem[ 6681] = 0;
disk_mem[ 6682] = 0;
disk_mem[ 6683] = 0;
disk_mem[ 6684] = 0;
disk_mem[ 6685] = 0;
disk_mem[ 6686] = 0;
disk_mem[ 6687] = 0;
disk_mem[ 6688] = 0;
disk_mem[ 6689] = 0;
disk_mem[ 6690] = 0;
disk_mem[ 6691] = 0;
disk_mem[ 6692] = 0;
disk_mem[ 6693] = 0;
disk_mem[ 6694] = 0;
disk_mem[ 6695] = 0;
disk_mem[ 6696] = 0;
disk_mem[ 6697] = 0;
disk_mem[ 6698] = 0;
disk_mem[ 6699] = 0;
disk_mem[ 6700] = 0;
disk_mem[ 6701] = 0;
disk_mem[ 6702] = 0;
disk_mem[ 6703] = 0;
disk_mem[ 6704] = 0;
disk_mem[ 6705] = 0;
disk_mem[ 6706] = 0;
disk_mem[ 6707] = 0;
disk_mem[ 6708] = 0;
disk_mem[ 6709] = 0;
disk_mem[ 6710] = 0;
disk_mem[ 6711] = 0;
disk_mem[ 6712] = 0;
disk_mem[ 6713] = 0;
disk_mem[ 6714] = 0;
disk_mem[ 6715] = 0;
disk_mem[ 6716] = 0;
disk_mem[ 6717] = 0;
disk_mem[ 6718] = 0;
disk_mem[ 6719] = 0;
disk_mem[ 6720] = 0;
disk_mem[ 6721] = 0;
disk_mem[ 6722] = 0;
disk_mem[ 6723] = 0;
disk_mem[ 6724] = 0;
disk_mem[ 6725] = 0;
disk_mem[ 6726] = 0;
disk_mem[ 6727] = 0;
disk_mem[ 6728] = 0;
disk_mem[ 6729] = 0;
disk_mem[ 6730] = 0;
disk_mem[ 6731] = 0;
disk_mem[ 6732] = 0;
disk_mem[ 6733] = 0;
disk_mem[ 6734] = 0;
disk_mem[ 6735] = 0;
disk_mem[ 6736] = 0;
disk_mem[ 6737] = 0;
disk_mem[ 6738] = 0;
disk_mem[ 6739] = 0;
disk_mem[ 6740] = 0;
disk_mem[ 6741] = 0;
disk_mem[ 6742] = 0;
disk_mem[ 6743] = 0;
disk_mem[ 6744] = 0;
disk_mem[ 6745] = 0;
disk_mem[ 6746] = 0;
disk_mem[ 6747] = 0;
disk_mem[ 6748] = 0;
disk_mem[ 6749] = 0;
disk_mem[ 6750] = 0;
disk_mem[ 6751] = 0;
disk_mem[ 6752] = 0;
disk_mem[ 6753] = 0;
disk_mem[ 6754] = 0;
disk_mem[ 6755] = 0;
disk_mem[ 6756] = 0;
disk_mem[ 6757] = 0;
disk_mem[ 6758] = 0;
disk_mem[ 6759] = 0;
disk_mem[ 6760] = 0;
disk_mem[ 6761] = 0;
disk_mem[ 6762] = 0;
disk_mem[ 6763] = 0;
disk_mem[ 6764] = 0;
disk_mem[ 6765] = 0;
disk_mem[ 6766] = 0;
disk_mem[ 6767] = 0;
disk_mem[ 6768] = 0;
disk_mem[ 6769] = 0;
disk_mem[ 6770] = 0;
disk_mem[ 6771] = 0;
disk_mem[ 6772] = 0;
disk_mem[ 6773] = 0;
disk_mem[ 6774] = 0;
disk_mem[ 6775] = 0;
disk_mem[ 6776] = 0;
disk_mem[ 6777] = 0;
disk_mem[ 6778] = 0;
disk_mem[ 6779] = 0;
disk_mem[ 6780] = 0;
disk_mem[ 6781] = 0;
disk_mem[ 6782] = 0;
disk_mem[ 6783] = 0;
disk_mem[ 6784] = 0;
disk_mem[ 6785] = 0;
disk_mem[ 6786] = 0;
disk_mem[ 6787] = 0;
disk_mem[ 6788] = 0;
disk_mem[ 6789] = 0;
disk_mem[ 6790] = 0;
disk_mem[ 6791] = 0;
disk_mem[ 6792] = 0;
disk_mem[ 6793] = 0;
disk_mem[ 6794] = 0;
disk_mem[ 6795] = 0;
disk_mem[ 6796] = 0;
disk_mem[ 6797] = 0;
disk_mem[ 6798] = 0;
disk_mem[ 6799] = 0;
disk_mem[ 6800] = 0;
disk_mem[ 6801] = 0;
disk_mem[ 6802] = 0;
disk_mem[ 6803] = 0;
disk_mem[ 6804] = 0;
disk_mem[ 6805] = 0;
disk_mem[ 6806] = 0;
disk_mem[ 6807] = 0;
disk_mem[ 6808] = 0;
disk_mem[ 6809] = 0;
disk_mem[ 6810] = 0;
disk_mem[ 6811] = 0;
disk_mem[ 6812] = 0;
disk_mem[ 6813] = 0;
disk_mem[ 6814] = 0;
disk_mem[ 6815] = 0;
disk_mem[ 6816] = 0;
disk_mem[ 6817] = 0;
disk_mem[ 6818] = 0;
disk_mem[ 6819] = 0;
disk_mem[ 6820] = 0;
disk_mem[ 6821] = 0;
disk_mem[ 6822] = 0;
disk_mem[ 6823] = 0;
disk_mem[ 6824] = 0;
disk_mem[ 6825] = 0;
disk_mem[ 6826] = 0;
disk_mem[ 6827] = 0;
disk_mem[ 6828] = 0;
disk_mem[ 6829] = 0;
disk_mem[ 6830] = 0;
disk_mem[ 6831] = 0;
disk_mem[ 6832] = 0;
disk_mem[ 6833] = 0;
disk_mem[ 6834] = 0;
disk_mem[ 6835] = 0;
disk_mem[ 6836] = 0;
disk_mem[ 6837] = 0;
disk_mem[ 6838] = 0;
disk_mem[ 6839] = 0;
disk_mem[ 6840] = 0;
disk_mem[ 6841] = 0;
disk_mem[ 6842] = 0;
disk_mem[ 6843] = 0;
disk_mem[ 6844] = 0;
disk_mem[ 6845] = 0;
disk_mem[ 6846] = 0;
disk_mem[ 6847] = 0;
disk_mem[ 6848] = 0;
disk_mem[ 6849] = 0;
disk_mem[ 6850] = 0;
disk_mem[ 6851] = 0;
disk_mem[ 6852] = 0;
disk_mem[ 6853] = 0;
disk_mem[ 6854] = 0;
disk_mem[ 6855] = 0;
disk_mem[ 6856] = 0;
disk_mem[ 6857] = 0;
disk_mem[ 6858] = 0;
disk_mem[ 6859] = 0;
disk_mem[ 6860] = 0;
disk_mem[ 6861] = 0;
disk_mem[ 6862] = 0;
disk_mem[ 6863] = 0;
disk_mem[ 6864] = 0;
disk_mem[ 6865] = 0;
disk_mem[ 6866] = 0;
disk_mem[ 6867] = 0;
disk_mem[ 6868] = 0;
disk_mem[ 6869] = 0;
disk_mem[ 6870] = 0;
disk_mem[ 6871] = 0;
disk_mem[ 6872] = 0;
disk_mem[ 6873] = 0;
disk_mem[ 6874] = 0;
disk_mem[ 6875] = 0;
disk_mem[ 6876] = 0;
disk_mem[ 6877] = 0;
disk_mem[ 6878] = 0;
disk_mem[ 6879] = 0;
disk_mem[ 6880] = 0;
disk_mem[ 6881] = 0;
disk_mem[ 6882] = 0;
disk_mem[ 6883] = 0;
disk_mem[ 6884] = 0;
disk_mem[ 6885] = 0;
disk_mem[ 6886] = 0;
disk_mem[ 6887] = 0;
disk_mem[ 6888] = 0;
disk_mem[ 6889] = 0;
disk_mem[ 6890] = 0;
disk_mem[ 6891] = 0;
disk_mem[ 6892] = 0;
disk_mem[ 6893] = 0;
disk_mem[ 6894] = 0;
disk_mem[ 6895] = 0;
disk_mem[ 6896] = 0;
disk_mem[ 6897] = 0;
disk_mem[ 6898] = 0;
disk_mem[ 6899] = 0;
disk_mem[ 6900] = 0;
disk_mem[ 6901] = 0;
disk_mem[ 6902] = 0;
disk_mem[ 6903] = 0;
disk_mem[ 6904] = 0;
disk_mem[ 6905] = 0;
disk_mem[ 6906] = 0;
disk_mem[ 6907] = 0;
disk_mem[ 6908] = 0;
disk_mem[ 6909] = 0;
disk_mem[ 6910] = 0;
disk_mem[ 6911] = 0;
disk_mem[ 6912] = 0;
disk_mem[ 6913] = 0;
disk_mem[ 6914] = 0;
disk_mem[ 6915] = 0;
disk_mem[ 6916] = 0;
disk_mem[ 6917] = 0;
disk_mem[ 6918] = 0;
disk_mem[ 6919] = 0;
disk_mem[ 6920] = 0;
disk_mem[ 6921] = 0;
disk_mem[ 6922] = 0;
disk_mem[ 6923] = 0;
disk_mem[ 6924] = 0;
disk_mem[ 6925] = 0;
disk_mem[ 6926] = 0;
disk_mem[ 6927] = 0;
disk_mem[ 6928] = 0;
disk_mem[ 6929] = 0;
disk_mem[ 6930] = 0;
disk_mem[ 6931] = 0;
disk_mem[ 6932] = 0;
disk_mem[ 6933] = 0;
disk_mem[ 6934] = 0;
disk_mem[ 6935] = 0;
disk_mem[ 6936] = 0;
disk_mem[ 6937] = 0;
disk_mem[ 6938] = 0;
disk_mem[ 6939] = 0;
disk_mem[ 6940] = 0;
disk_mem[ 6941] = 0;
disk_mem[ 6942] = 0;
disk_mem[ 6943] = 0;
disk_mem[ 6944] = 0;
disk_mem[ 6945] = 0;
disk_mem[ 6946] = 0;
disk_mem[ 6947] = 0;
disk_mem[ 6948] = 0;
disk_mem[ 6949] = 0;
disk_mem[ 6950] = 0;
disk_mem[ 6951] = 0;
disk_mem[ 6952] = 0;
disk_mem[ 6953] = 0;
disk_mem[ 6954] = 0;
disk_mem[ 6955] = 0;
disk_mem[ 6956] = 0;
disk_mem[ 6957] = 0;
disk_mem[ 6958] = 0;
disk_mem[ 6959] = 0;
disk_mem[ 6960] = 0;
disk_mem[ 6961] = 0;
disk_mem[ 6962] = 0;
disk_mem[ 6963] = 0;
disk_mem[ 6964] = 0;
disk_mem[ 6965] = 0;
disk_mem[ 6966] = 0;
disk_mem[ 6967] = 0;
disk_mem[ 6968] = 0;
disk_mem[ 6969] = 0;
disk_mem[ 6970] = 0;
disk_mem[ 6971] = 0;
disk_mem[ 6972] = 0;
disk_mem[ 6973] = 0;
disk_mem[ 6974] = 0;
disk_mem[ 6975] = 0;
disk_mem[ 6976] = 0;
disk_mem[ 6977] = 0;
disk_mem[ 6978] = 0;
disk_mem[ 6979] = 0;
disk_mem[ 6980] = 0;
disk_mem[ 6981] = 0;
disk_mem[ 6982] = 0;
disk_mem[ 6983] = 0;
disk_mem[ 6984] = 0;
disk_mem[ 6985] = 0;
disk_mem[ 6986] = 0;
disk_mem[ 6987] = 0;
disk_mem[ 6988] = 0;
disk_mem[ 6989] = 0;
disk_mem[ 6990] = 0;
disk_mem[ 6991] = 0;
disk_mem[ 6992] = 0;
disk_mem[ 6993] = 0;
disk_mem[ 6994] = 0;
disk_mem[ 6995] = 0;
disk_mem[ 6996] = 0;
disk_mem[ 6997] = 0;
disk_mem[ 6998] = 0;
disk_mem[ 6999] = 0;
disk_mem[ 7000] = 0;
disk_mem[ 7001] = 0;
disk_mem[ 7002] = 0;
disk_mem[ 7003] = 0;
disk_mem[ 7004] = 0;
disk_mem[ 7005] = 0;
disk_mem[ 7006] = 0;
disk_mem[ 7007] = 0;
disk_mem[ 7008] = 0;
disk_mem[ 7009] = 0;
disk_mem[ 7010] = 0;
disk_mem[ 7011] = 0;
disk_mem[ 7012] = 0;
disk_mem[ 7013] = 0;
disk_mem[ 7014] = 0;
disk_mem[ 7015] = 0;
disk_mem[ 7016] = 0;
disk_mem[ 7017] = 0;
disk_mem[ 7018] = 0;
disk_mem[ 7019] = 0;
disk_mem[ 7020] = 0;
disk_mem[ 7021] = 0;
disk_mem[ 7022] = 0;
disk_mem[ 7023] = 0;
disk_mem[ 7024] = 0;
disk_mem[ 7025] = 0;
disk_mem[ 7026] = 0;
disk_mem[ 7027] = 0;
disk_mem[ 7028] = 0;
disk_mem[ 7029] = 0;
disk_mem[ 7030] = 0;
disk_mem[ 7031] = 0;
disk_mem[ 7032] = 0;
disk_mem[ 7033] = 0;
disk_mem[ 7034] = 0;
disk_mem[ 7035] = 0;
disk_mem[ 7036] = 0;
disk_mem[ 7037] = 0;
disk_mem[ 7038] = 0;
disk_mem[ 7039] = 0;
disk_mem[ 7040] = 0;
disk_mem[ 7041] = 0;
disk_mem[ 7042] = 0;
disk_mem[ 7043] = 0;
disk_mem[ 7044] = 0;
disk_mem[ 7045] = 0;
disk_mem[ 7046] = 0;
disk_mem[ 7047] = 0;
disk_mem[ 7048] = 0;
disk_mem[ 7049] = 0;
disk_mem[ 7050] = 0;
disk_mem[ 7051] = 0;
disk_mem[ 7052] = 0;
disk_mem[ 7053] = 0;
disk_mem[ 7054] = 0;
disk_mem[ 7055] = 0;
disk_mem[ 7056] = 0;
disk_mem[ 7057] = 0;
disk_mem[ 7058] = 0;
disk_mem[ 7059] = 0;
disk_mem[ 7060] = 0;
disk_mem[ 7061] = 0;
disk_mem[ 7062] = 0;
disk_mem[ 7063] = 0;
disk_mem[ 7064] = 0;
disk_mem[ 7065] = 0;
disk_mem[ 7066] = 0;
disk_mem[ 7067] = 0;
disk_mem[ 7068] = 0;
disk_mem[ 7069] = 0;
disk_mem[ 7070] = 0;
disk_mem[ 7071] = 0;
disk_mem[ 7072] = 0;
disk_mem[ 7073] = 0;
disk_mem[ 7074] = 0;
disk_mem[ 7075] = 0;
disk_mem[ 7076] = 0;
disk_mem[ 7077] = 0;
disk_mem[ 7078] = 0;
disk_mem[ 7079] = 0;
disk_mem[ 7080] = 0;
disk_mem[ 7081] = 0;
disk_mem[ 7082] = 0;
disk_mem[ 7083] = 0;
disk_mem[ 7084] = 0;
disk_mem[ 7085] = 0;
disk_mem[ 7086] = 0;
disk_mem[ 7087] = 0;
disk_mem[ 7088] = 0;
disk_mem[ 7089] = 0;
disk_mem[ 7090] = 0;
disk_mem[ 7091] = 0;
disk_mem[ 7092] = 0;
disk_mem[ 7093] = 0;
disk_mem[ 7094] = 0;
disk_mem[ 7095] = 0;
disk_mem[ 7096] = 0;
disk_mem[ 7097] = 0;
disk_mem[ 7098] = 0;
disk_mem[ 7099] = 0;
disk_mem[ 7100] = 0;
disk_mem[ 7101] = 0;
disk_mem[ 7102] = 0;
disk_mem[ 7103] = 0;
disk_mem[ 7104] = 0;
disk_mem[ 7105] = 0;
disk_mem[ 7106] = 0;
disk_mem[ 7107] = 0;
disk_mem[ 7108] = 0;
disk_mem[ 7109] = 0;
disk_mem[ 7110] = 0;
disk_mem[ 7111] = 0;
disk_mem[ 7112] = 0;
disk_mem[ 7113] = 0;
disk_mem[ 7114] = 0;
disk_mem[ 7115] = 0;
disk_mem[ 7116] = 0;
disk_mem[ 7117] = 0;
disk_mem[ 7118] = 0;
disk_mem[ 7119] = 0;
disk_mem[ 7120] = 0;
disk_mem[ 7121] = 0;
disk_mem[ 7122] = 0;
disk_mem[ 7123] = 0;
disk_mem[ 7124] = 0;
disk_mem[ 7125] = 0;
disk_mem[ 7126] = 0;
disk_mem[ 7127] = 0;
disk_mem[ 7128] = 0;
disk_mem[ 7129] = 0;
disk_mem[ 7130] = 0;
disk_mem[ 7131] = 0;
disk_mem[ 7132] = 0;
disk_mem[ 7133] = 0;
disk_mem[ 7134] = 0;
disk_mem[ 7135] = 0;
disk_mem[ 7136] = 0;
disk_mem[ 7137] = 0;
disk_mem[ 7138] = 0;
disk_mem[ 7139] = 0;
disk_mem[ 7140] = 0;
disk_mem[ 7141] = 0;
disk_mem[ 7142] = 0;
disk_mem[ 7143] = 0;
disk_mem[ 7144] = 0;
disk_mem[ 7145] = 0;
disk_mem[ 7146] = 0;
disk_mem[ 7147] = 0;
disk_mem[ 7148] = 0;
disk_mem[ 7149] = 0;
disk_mem[ 7150] = 0;
disk_mem[ 7151] = 0;
disk_mem[ 7152] = 0;
disk_mem[ 7153] = 0;
disk_mem[ 7154] = 0;
disk_mem[ 7155] = 0;
disk_mem[ 7156] = 0;
disk_mem[ 7157] = 0;
disk_mem[ 7158] = 0;
disk_mem[ 7159] = 0;
disk_mem[ 7160] = 0;
disk_mem[ 7161] = 0;
disk_mem[ 7162] = 0;
disk_mem[ 7163] = 0;
disk_mem[ 7164] = 0;
disk_mem[ 7165] = 0;
disk_mem[ 7166] = 0;
disk_mem[ 7167] = 0;
disk_mem[ 7168] = 0;
disk_mem[ 7169] = 0;
disk_mem[ 7170] = 0;
disk_mem[ 7171] = 0;
disk_mem[ 7172] = 0;
disk_mem[ 7173] = 0;
disk_mem[ 7174] = 0;
disk_mem[ 7175] = 0;
disk_mem[ 7176] = 0;
disk_mem[ 7177] = 0;
disk_mem[ 7178] = 0;
disk_mem[ 7179] = 0;
disk_mem[ 7180] = 0;
disk_mem[ 7181] = 0;
disk_mem[ 7182] = 0;
disk_mem[ 7183] = 0;
disk_mem[ 7184] = 0;
disk_mem[ 7185] = 0;
disk_mem[ 7186] = 0;
disk_mem[ 7187] = 0;
disk_mem[ 7188] = 0;
disk_mem[ 7189] = 0;
disk_mem[ 7190] = 0;
disk_mem[ 7191] = 0;
disk_mem[ 7192] = 0;
disk_mem[ 7193] = 0;
disk_mem[ 7194] = 0;
disk_mem[ 7195] = 0;
disk_mem[ 7196] = 0;
disk_mem[ 7197] = 0;
disk_mem[ 7198] = 0;
disk_mem[ 7199] = 0;
disk_mem[ 7200] = 0;
disk_mem[ 7201] = 0;
disk_mem[ 7202] = 0;
disk_mem[ 7203] = 0;
disk_mem[ 7204] = 0;
disk_mem[ 7205] = 0;
disk_mem[ 7206] = 0;
disk_mem[ 7207] = 0;
disk_mem[ 7208] = 0;
disk_mem[ 7209] = 0;
disk_mem[ 7210] = 0;
disk_mem[ 7211] = 0;
disk_mem[ 7212] = 0;
disk_mem[ 7213] = 0;
disk_mem[ 7214] = 0;
disk_mem[ 7215] = 0;
disk_mem[ 7216] = 0;
disk_mem[ 7217] = 0;
disk_mem[ 7218] = 0;
disk_mem[ 7219] = 0;
disk_mem[ 7220] = 0;
disk_mem[ 7221] = 0;
disk_mem[ 7222] = 0;
disk_mem[ 7223] = 0;
disk_mem[ 7224] = 0;
disk_mem[ 7225] = 0;
disk_mem[ 7226] = 0;
disk_mem[ 7227] = 0;
disk_mem[ 7228] = 0;
disk_mem[ 7229] = 0;
disk_mem[ 7230] = 0;
disk_mem[ 7231] = 0;
disk_mem[ 7232] = 0;
disk_mem[ 7233] = 0;
disk_mem[ 7234] = 0;
disk_mem[ 7235] = 0;
disk_mem[ 7236] = 0;
disk_mem[ 7237] = 0;
disk_mem[ 7238] = 0;
disk_mem[ 7239] = 0;
disk_mem[ 7240] = 0;
disk_mem[ 7241] = 0;
disk_mem[ 7242] = 0;
disk_mem[ 7243] = 0;
disk_mem[ 7244] = 0;
disk_mem[ 7245] = 0;
disk_mem[ 7246] = 0;
disk_mem[ 7247] = 0;
disk_mem[ 7248] = 0;
disk_mem[ 7249] = 0;
disk_mem[ 7250] = 0;
disk_mem[ 7251] = 0;
disk_mem[ 7252] = 0;
disk_mem[ 7253] = 0;
disk_mem[ 7254] = 0;
disk_mem[ 7255] = 0;
disk_mem[ 7256] = 0;
disk_mem[ 7257] = 0;
disk_mem[ 7258] = 0;
disk_mem[ 7259] = 0;
disk_mem[ 7260] = 0;
disk_mem[ 7261] = 0;
disk_mem[ 7262] = 0;
disk_mem[ 7263] = 0;
disk_mem[ 7264] = 0;
disk_mem[ 7265] = 0;
disk_mem[ 7266] = 0;
disk_mem[ 7267] = 0;
disk_mem[ 7268] = 0;
disk_mem[ 7269] = 0;
disk_mem[ 7270] = 0;
disk_mem[ 7271] = 0;
disk_mem[ 7272] = 0;
disk_mem[ 7273] = 0;
disk_mem[ 7274] = 0;
disk_mem[ 7275] = 0;
disk_mem[ 7276] = 0;
disk_mem[ 7277] = 0;
disk_mem[ 7278] = 0;
disk_mem[ 7279] = 0;
disk_mem[ 7280] = 0;
disk_mem[ 7281] = 0;
disk_mem[ 7282] = 0;
disk_mem[ 7283] = 0;
disk_mem[ 7284] = 0;
disk_mem[ 7285] = 0;
disk_mem[ 7286] = 0;
disk_mem[ 7287] = 0;
disk_mem[ 7288] = 0;
disk_mem[ 7289] = 0;
disk_mem[ 7290] = 0;
disk_mem[ 7291] = 0;
disk_mem[ 7292] = 0;
disk_mem[ 7293] = 0;
disk_mem[ 7294] = 0;
disk_mem[ 7295] = 0;
disk_mem[ 7296] = 0;
disk_mem[ 7297] = 0;
disk_mem[ 7298] = 0;
disk_mem[ 7299] = 0;
disk_mem[ 7300] = 0;
disk_mem[ 7301] = 0;
disk_mem[ 7302] = 0;
disk_mem[ 7303] = 0;
disk_mem[ 7304] = 0;
disk_mem[ 7305] = 0;
disk_mem[ 7306] = 0;
disk_mem[ 7307] = 0;
disk_mem[ 7308] = 0;
disk_mem[ 7309] = 0;
disk_mem[ 7310] = 0;
disk_mem[ 7311] = 0;
disk_mem[ 7312] = 0;
disk_mem[ 7313] = 0;
disk_mem[ 7314] = 0;
disk_mem[ 7315] = 0;
disk_mem[ 7316] = 0;
disk_mem[ 7317] = 0;
disk_mem[ 7318] = 0;
disk_mem[ 7319] = 0;
disk_mem[ 7320] = 0;
disk_mem[ 7321] = 0;
disk_mem[ 7322] = 0;
disk_mem[ 7323] = 0;
disk_mem[ 7324] = 0;
disk_mem[ 7325] = 0;
disk_mem[ 7326] = 0;
disk_mem[ 7327] = 0;
disk_mem[ 7328] = 0;
disk_mem[ 7329] = 0;
disk_mem[ 7330] = 0;
disk_mem[ 7331] = 0;
disk_mem[ 7332] = 0;
disk_mem[ 7333] = 0;
disk_mem[ 7334] = 0;
disk_mem[ 7335] = 0;
disk_mem[ 7336] = 0;
disk_mem[ 7337] = 0;
disk_mem[ 7338] = 0;
disk_mem[ 7339] = 0;
disk_mem[ 7340] = 0;
disk_mem[ 7341] = 0;
disk_mem[ 7342] = 0;
disk_mem[ 7343] = 0;
disk_mem[ 7344] = 0;
disk_mem[ 7345] = 0;
disk_mem[ 7346] = 0;
disk_mem[ 7347] = 0;
disk_mem[ 7348] = 0;
disk_mem[ 7349] = 0;
disk_mem[ 7350] = 0;
disk_mem[ 7351] = 0;
disk_mem[ 7352] = 0;
disk_mem[ 7353] = 0;
disk_mem[ 7354] = 0;
disk_mem[ 7355] = 0;
disk_mem[ 7356] = 0;
disk_mem[ 7357] = 0;
disk_mem[ 7358] = 0;
disk_mem[ 7359] = 0;
disk_mem[ 7360] = 0;
disk_mem[ 7361] = 0;
disk_mem[ 7362] = 0;
disk_mem[ 7363] = 0;
disk_mem[ 7364] = 0;
disk_mem[ 7365] = 0;
disk_mem[ 7366] = 0;
disk_mem[ 7367] = 0;
disk_mem[ 7368] = 0;
disk_mem[ 7369] = 0;
disk_mem[ 7370] = 0;
disk_mem[ 7371] = 0;
disk_mem[ 7372] = 0;
disk_mem[ 7373] = 0;
disk_mem[ 7374] = 0;
disk_mem[ 7375] = 0;
disk_mem[ 7376] = 0;
disk_mem[ 7377] = 0;
disk_mem[ 7378] = 0;
disk_mem[ 7379] = 0;
disk_mem[ 7380] = 0;
disk_mem[ 7381] = 0;
disk_mem[ 7382] = 0;
disk_mem[ 7383] = 0;
disk_mem[ 7384] = 0;
disk_mem[ 7385] = 0;
disk_mem[ 7386] = 0;
disk_mem[ 7387] = 0;
disk_mem[ 7388] = 0;
disk_mem[ 7389] = 0;
disk_mem[ 7390] = 0;
disk_mem[ 7391] = 0;
disk_mem[ 7392] = 0;
disk_mem[ 7393] = 0;
disk_mem[ 7394] = 0;
disk_mem[ 7395] = 0;
disk_mem[ 7396] = 0;
disk_mem[ 7397] = 0;
disk_mem[ 7398] = 0;
disk_mem[ 7399] = 0;
disk_mem[ 7400] = 0;
disk_mem[ 7401] = 0;
disk_mem[ 7402] = 0;
disk_mem[ 7403] = 0;
disk_mem[ 7404] = 0;
disk_mem[ 7405] = 0;
disk_mem[ 7406] = 0;
disk_mem[ 7407] = 0;
disk_mem[ 7408] = 0;
disk_mem[ 7409] = 0;
disk_mem[ 7410] = 0;
disk_mem[ 7411] = 0;
disk_mem[ 7412] = 0;
disk_mem[ 7413] = 0;
disk_mem[ 7414] = 0;
disk_mem[ 7415] = 0;
disk_mem[ 7416] = 0;
disk_mem[ 7417] = 0;
disk_mem[ 7418] = 0;
disk_mem[ 7419] = 0;
disk_mem[ 7420] = 0;
disk_mem[ 7421] = 0;
disk_mem[ 7422] = 0;
disk_mem[ 7423] = 0;
disk_mem[ 7424] = 0;
disk_mem[ 7425] = 0;
disk_mem[ 7426] = 0;
disk_mem[ 7427] = 0;
disk_mem[ 7428] = 0;
disk_mem[ 7429] = 0;
disk_mem[ 7430] = 0;
disk_mem[ 7431] = 0;
disk_mem[ 7432] = 0;
disk_mem[ 7433] = 0;
disk_mem[ 7434] = 0;
disk_mem[ 7435] = 0;
disk_mem[ 7436] = 0;
disk_mem[ 7437] = 0;
disk_mem[ 7438] = 0;
disk_mem[ 7439] = 0;
disk_mem[ 7440] = 0;
disk_mem[ 7441] = 0;
disk_mem[ 7442] = 0;
disk_mem[ 7443] = 0;
disk_mem[ 7444] = 0;
disk_mem[ 7445] = 0;
disk_mem[ 7446] = 0;
disk_mem[ 7447] = 0;
disk_mem[ 7448] = 0;
disk_mem[ 7449] = 0;
disk_mem[ 7450] = 0;
disk_mem[ 7451] = 0;
disk_mem[ 7452] = 0;
disk_mem[ 7453] = 0;
disk_mem[ 7454] = 0;
disk_mem[ 7455] = 0;
disk_mem[ 7456] = 0;
disk_mem[ 7457] = 0;
disk_mem[ 7458] = 0;
disk_mem[ 7459] = 0;
disk_mem[ 7460] = 0;
disk_mem[ 7461] = 0;
disk_mem[ 7462] = 0;
disk_mem[ 7463] = 0;
disk_mem[ 7464] = 0;
disk_mem[ 7465] = 0;
disk_mem[ 7466] = 0;
disk_mem[ 7467] = 0;
disk_mem[ 7468] = 0;
disk_mem[ 7469] = 0;
disk_mem[ 7470] = 0;
disk_mem[ 7471] = 0;
disk_mem[ 7472] = 0;
disk_mem[ 7473] = 0;
disk_mem[ 7474] = 0;
disk_mem[ 7475] = 0;
disk_mem[ 7476] = 0;
disk_mem[ 7477] = 0;
disk_mem[ 7478] = 0;
disk_mem[ 7479] = 0;
disk_mem[ 7480] = 0;
disk_mem[ 7481] = 0;
disk_mem[ 7482] = 0;
disk_mem[ 7483] = 0;
disk_mem[ 7484] = 0;
disk_mem[ 7485] = 0;
disk_mem[ 7486] = 0;
disk_mem[ 7487] = 0;
disk_mem[ 7488] = 0;
disk_mem[ 7489] = 0;
disk_mem[ 7490] = 0;
disk_mem[ 7491] = 0;
disk_mem[ 7492] = 0;
disk_mem[ 7493] = 0;
disk_mem[ 7494] = 0;
disk_mem[ 7495] = 0;
disk_mem[ 7496] = 0;
disk_mem[ 7497] = 0;
disk_mem[ 7498] = 0;
disk_mem[ 7499] = 0;
disk_mem[ 7500] = 0;
disk_mem[ 7501] = 0;
disk_mem[ 7502] = 0;
disk_mem[ 7503] = 0;
disk_mem[ 7504] = 0;
disk_mem[ 7505] = 0;
disk_mem[ 7506] = 0;
disk_mem[ 7507] = 0;
disk_mem[ 7508] = 0;
disk_mem[ 7509] = 0;
disk_mem[ 7510] = 0;
disk_mem[ 7511] = 0;
disk_mem[ 7512] = 0;
disk_mem[ 7513] = 0;
disk_mem[ 7514] = 0;
disk_mem[ 7515] = 0;
disk_mem[ 7516] = 0;
disk_mem[ 7517] = 0;
disk_mem[ 7518] = 0;
disk_mem[ 7519] = 0;
disk_mem[ 7520] = 0;
disk_mem[ 7521] = 0;
disk_mem[ 7522] = 0;
disk_mem[ 7523] = 0;
disk_mem[ 7524] = 0;
disk_mem[ 7525] = 0;
disk_mem[ 7526] = 0;
disk_mem[ 7527] = 0;
disk_mem[ 7528] = 0;
disk_mem[ 7529] = 0;
disk_mem[ 7530] = 0;
disk_mem[ 7531] = 0;
disk_mem[ 7532] = 0;
disk_mem[ 7533] = 0;
disk_mem[ 7534] = 0;
disk_mem[ 7535] = 0;
disk_mem[ 7536] = 0;
disk_mem[ 7537] = 0;
disk_mem[ 7538] = 0;
disk_mem[ 7539] = 0;
disk_mem[ 7540] = 0;
disk_mem[ 7541] = 0;
disk_mem[ 7542] = 0;
disk_mem[ 7543] = 0;
disk_mem[ 7544] = 0;
disk_mem[ 7545] = 0;
disk_mem[ 7546] = 0;
disk_mem[ 7547] = 0;
disk_mem[ 7548] = 0;
disk_mem[ 7549] = 0;
disk_mem[ 7550] = 0;
disk_mem[ 7551] = 0;
disk_mem[ 7552] = 0;
disk_mem[ 7553] = 0;
disk_mem[ 7554] = 0;
disk_mem[ 7555] = 0;
disk_mem[ 7556] = 0;
disk_mem[ 7557] = 0;
disk_mem[ 7558] = 0;
disk_mem[ 7559] = 0;
disk_mem[ 7560] = 0;
disk_mem[ 7561] = 0;
disk_mem[ 7562] = 0;
disk_mem[ 7563] = 0;
disk_mem[ 7564] = 0;
disk_mem[ 7565] = 0;
disk_mem[ 7566] = 0;
disk_mem[ 7567] = 0;
disk_mem[ 7568] = 0;
disk_mem[ 7569] = 0;
disk_mem[ 7570] = 0;
disk_mem[ 7571] = 0;
disk_mem[ 7572] = 0;
disk_mem[ 7573] = 0;
disk_mem[ 7574] = 0;
disk_mem[ 7575] = 0;
disk_mem[ 7576] = 0;
disk_mem[ 7577] = 0;
disk_mem[ 7578] = 0;
disk_mem[ 7579] = 0;
disk_mem[ 7580] = 0;
disk_mem[ 7581] = 0;
disk_mem[ 7582] = 0;
disk_mem[ 7583] = 0;
disk_mem[ 7584] = 0;
disk_mem[ 7585] = 0;
disk_mem[ 7586] = 0;
disk_mem[ 7587] = 0;
disk_mem[ 7588] = 0;
disk_mem[ 7589] = 0;
disk_mem[ 7590] = 0;
disk_mem[ 7591] = 0;
disk_mem[ 7592] = 0;
disk_mem[ 7593] = 0;
disk_mem[ 7594] = 0;
disk_mem[ 7595] = 0;
disk_mem[ 7596] = 0;
disk_mem[ 7597] = 0;
disk_mem[ 7598] = 0;
disk_mem[ 7599] = 0;
disk_mem[ 7600] = 0;
disk_mem[ 7601] = 0;
disk_mem[ 7602] = 0;
disk_mem[ 7603] = 0;
disk_mem[ 7604] = 0;
disk_mem[ 7605] = 0;
disk_mem[ 7606] = 0;
disk_mem[ 7607] = 0;
disk_mem[ 7608] = 0;
disk_mem[ 7609] = 0;
disk_mem[ 7610] = 0;
disk_mem[ 7611] = 0;
disk_mem[ 7612] = 0;
disk_mem[ 7613] = 0;
disk_mem[ 7614] = 0;
disk_mem[ 7615] = 0;
disk_mem[ 7616] = 0;
disk_mem[ 7617] = 0;
disk_mem[ 7618] = 0;
disk_mem[ 7619] = 0;
disk_mem[ 7620] = 0;
disk_mem[ 7621] = 0;
disk_mem[ 7622] = 0;
disk_mem[ 7623] = 0;
disk_mem[ 7624] = 0;
disk_mem[ 7625] = 0;
disk_mem[ 7626] = 0;
disk_mem[ 7627] = 0;
disk_mem[ 7628] = 0;
disk_mem[ 7629] = 0;
disk_mem[ 7630] = 0;
disk_mem[ 7631] = 0;
disk_mem[ 7632] = 0;
disk_mem[ 7633] = 0;
disk_mem[ 7634] = 0;
disk_mem[ 7635] = 0;
disk_mem[ 7636] = 0;
disk_mem[ 7637] = 0;
disk_mem[ 7638] = 0;
disk_mem[ 7639] = 0;
disk_mem[ 7640] = 0;
disk_mem[ 7641] = 0;
disk_mem[ 7642] = 0;
disk_mem[ 7643] = 0;
disk_mem[ 7644] = 0;
disk_mem[ 7645] = 0;
disk_mem[ 7646] = 0;
disk_mem[ 7647] = 0;
disk_mem[ 7648] = 0;
disk_mem[ 7649] = 0;
disk_mem[ 7650] = 0;
disk_mem[ 7651] = 0;
disk_mem[ 7652] = 0;
disk_mem[ 7653] = 0;
disk_mem[ 7654] = 0;
disk_mem[ 7655] = 0;
disk_mem[ 7656] = 0;
disk_mem[ 7657] = 0;
disk_mem[ 7658] = 0;
disk_mem[ 7659] = 0;
disk_mem[ 7660] = 0;
disk_mem[ 7661] = 0;
disk_mem[ 7662] = 0;
disk_mem[ 7663] = 0;
disk_mem[ 7664] = 0;
disk_mem[ 7665] = 0;
disk_mem[ 7666] = 0;
disk_mem[ 7667] = 0;
disk_mem[ 7668] = 0;
disk_mem[ 7669] = 0;
disk_mem[ 7670] = 0;
disk_mem[ 7671] = 0;
disk_mem[ 7672] = 0;
disk_mem[ 7673] = 0;
disk_mem[ 7674] = 0;
disk_mem[ 7675] = 0;
disk_mem[ 7676] = 0;
disk_mem[ 7677] = 0;
disk_mem[ 7678] = 0;
disk_mem[ 7679] = 0;
disk_mem[ 7680] = 0;
disk_mem[ 7681] = 0;
disk_mem[ 7682] = 0;
disk_mem[ 7683] = 0;
disk_mem[ 7684] = 0;
disk_mem[ 7685] = 0;
disk_mem[ 7686] = 0;
disk_mem[ 7687] = 0;
disk_mem[ 7688] = 0;
disk_mem[ 7689] = 0;
disk_mem[ 7690] = 0;
disk_mem[ 7691] = 0;
disk_mem[ 7692] = 0;
disk_mem[ 7693] = 0;
disk_mem[ 7694] = 0;
disk_mem[ 7695] = 0;
disk_mem[ 7696] = 0;
disk_mem[ 7697] = 0;
disk_mem[ 7698] = 0;
disk_mem[ 7699] = 0;
disk_mem[ 7700] = 0;
disk_mem[ 7701] = 0;
disk_mem[ 7702] = 0;
disk_mem[ 7703] = 0;
disk_mem[ 7704] = 0;
disk_mem[ 7705] = 0;
disk_mem[ 7706] = 0;
disk_mem[ 7707] = 0;
disk_mem[ 7708] = 0;
disk_mem[ 7709] = 0;
disk_mem[ 7710] = 0;
disk_mem[ 7711] = 0;
disk_mem[ 7712] = 0;
disk_mem[ 7713] = 0;
disk_mem[ 7714] = 0;
disk_mem[ 7715] = 0;
disk_mem[ 7716] = 0;
disk_mem[ 7717] = 0;
disk_mem[ 7718] = 0;
disk_mem[ 7719] = 0;
disk_mem[ 7720] = 0;
disk_mem[ 7721] = 0;
disk_mem[ 7722] = 0;
disk_mem[ 7723] = 0;
disk_mem[ 7724] = 0;
disk_mem[ 7725] = 0;
disk_mem[ 7726] = 0;
disk_mem[ 7727] = 0;
disk_mem[ 7728] = 0;
disk_mem[ 7729] = 0;
disk_mem[ 7730] = 0;
disk_mem[ 7731] = 0;
disk_mem[ 7732] = 0;
disk_mem[ 7733] = 0;
disk_mem[ 7734] = 0;
disk_mem[ 7735] = 0;
disk_mem[ 7736] = 0;
disk_mem[ 7737] = 0;
disk_mem[ 7738] = 0;
disk_mem[ 7739] = 0;
disk_mem[ 7740] = 0;
disk_mem[ 7741] = 0;
disk_mem[ 7742] = 0;
disk_mem[ 7743] = 0;
disk_mem[ 7744] = 0;
disk_mem[ 7745] = 0;
disk_mem[ 7746] = 0;
disk_mem[ 7747] = 0;
disk_mem[ 7748] = 0;
disk_mem[ 7749] = 0;
disk_mem[ 7750] = 0;
disk_mem[ 7751] = 0;
disk_mem[ 7752] = 0;
disk_mem[ 7753] = 0;
disk_mem[ 7754] = 0;
disk_mem[ 7755] = 0;
disk_mem[ 7756] = 0;
disk_mem[ 7757] = 0;
disk_mem[ 7758] = 0;
disk_mem[ 7759] = 0;
disk_mem[ 7760] = 0;
disk_mem[ 7761] = 0;
disk_mem[ 7762] = 0;
disk_mem[ 7763] = 0;
disk_mem[ 7764] = 0;
disk_mem[ 7765] = 0;
disk_mem[ 7766] = 0;
disk_mem[ 7767] = 0;
disk_mem[ 7768] = 0;
disk_mem[ 7769] = 0;
disk_mem[ 7770] = 0;
disk_mem[ 7771] = 0;
disk_mem[ 7772] = 0;
disk_mem[ 7773] = 0;
disk_mem[ 7774] = 0;
disk_mem[ 7775] = 0;
disk_mem[ 7776] = 0;
disk_mem[ 7777] = 0;
disk_mem[ 7778] = 0;
disk_mem[ 7779] = 0;
disk_mem[ 7780] = 0;
disk_mem[ 7781] = 0;
disk_mem[ 7782] = 0;
disk_mem[ 7783] = 0;
disk_mem[ 7784] = 0;
disk_mem[ 7785] = 0;
disk_mem[ 7786] = 0;
disk_mem[ 7787] = 0;
disk_mem[ 7788] = 0;
disk_mem[ 7789] = 0;
disk_mem[ 7790] = 0;
disk_mem[ 7791] = 0;
disk_mem[ 7792] = 0;
disk_mem[ 7793] = 0;
disk_mem[ 7794] = 0;
disk_mem[ 7795] = 0;
disk_mem[ 7796] = 0;
disk_mem[ 7797] = 0;
disk_mem[ 7798] = 0;
disk_mem[ 7799] = 0;
disk_mem[ 7800] = 0;
disk_mem[ 7801] = 0;
disk_mem[ 7802] = 0;
disk_mem[ 7803] = 0;
disk_mem[ 7804] = 0;
disk_mem[ 7805] = 0;
disk_mem[ 7806] = 0;
disk_mem[ 7807] = 0;
disk_mem[ 7808] = 0;
disk_mem[ 7809] = 0;
disk_mem[ 7810] = 0;
disk_mem[ 7811] = 0;
disk_mem[ 7812] = 0;
disk_mem[ 7813] = 0;
disk_mem[ 7814] = 0;
disk_mem[ 7815] = 0;
disk_mem[ 7816] = 0;
disk_mem[ 7817] = 0;
disk_mem[ 7818] = 0;
disk_mem[ 7819] = 0;
disk_mem[ 7820] = 0;
disk_mem[ 7821] = 0;
disk_mem[ 7822] = 0;
disk_mem[ 7823] = 0;
disk_mem[ 7824] = 0;
disk_mem[ 7825] = 0;
disk_mem[ 7826] = 0;
disk_mem[ 7827] = 0;
disk_mem[ 7828] = 0;
disk_mem[ 7829] = 0;
disk_mem[ 7830] = 0;
disk_mem[ 7831] = 0;
disk_mem[ 7832] = 0;
disk_mem[ 7833] = 0;
disk_mem[ 7834] = 0;
disk_mem[ 7835] = 0;
disk_mem[ 7836] = 0;
disk_mem[ 7837] = 0;
disk_mem[ 7838] = 0;
disk_mem[ 7839] = 0;
disk_mem[ 7840] = 0;
disk_mem[ 7841] = 0;
disk_mem[ 7842] = 0;
disk_mem[ 7843] = 0;
disk_mem[ 7844] = 0;
disk_mem[ 7845] = 0;
disk_mem[ 7846] = 0;
disk_mem[ 7847] = 0;
disk_mem[ 7848] = 0;
disk_mem[ 7849] = 0;
disk_mem[ 7850] = 0;
disk_mem[ 7851] = 0;
disk_mem[ 7852] = 0;
disk_mem[ 7853] = 0;
disk_mem[ 7854] = 0;
disk_mem[ 7855] = 0;
disk_mem[ 7856] = 0;
disk_mem[ 7857] = 0;
disk_mem[ 7858] = 0;
disk_mem[ 7859] = 0;
disk_mem[ 7860] = 0;
disk_mem[ 7861] = 0;
disk_mem[ 7862] = 0;
disk_mem[ 7863] = 0;
disk_mem[ 7864] = 0;
disk_mem[ 7865] = 0;
disk_mem[ 7866] = 0;
disk_mem[ 7867] = 0;
disk_mem[ 7868] = 0;
disk_mem[ 7869] = 0;
disk_mem[ 7870] = 0;
disk_mem[ 7871] = 0;
disk_mem[ 7872] = 0;
disk_mem[ 7873] = 0;
disk_mem[ 7874] = 0;
disk_mem[ 7875] = 0;
disk_mem[ 7876] = 0;
disk_mem[ 7877] = 0;
disk_mem[ 7878] = 0;
disk_mem[ 7879] = 0;
disk_mem[ 7880] = 0;
disk_mem[ 7881] = 0;
disk_mem[ 7882] = 0;
disk_mem[ 7883] = 0;
disk_mem[ 7884] = 0;
disk_mem[ 7885] = 0;
disk_mem[ 7886] = 0;
disk_mem[ 7887] = 0;
disk_mem[ 7888] = 0;
disk_mem[ 7889] = 0;
disk_mem[ 7890] = 0;
disk_mem[ 7891] = 0;
disk_mem[ 7892] = 0;
disk_mem[ 7893] = 0;
disk_mem[ 7894] = 0;
disk_mem[ 7895] = 0;
disk_mem[ 7896] = 0;
disk_mem[ 7897] = 0;
disk_mem[ 7898] = 0;
disk_mem[ 7899] = 0;
disk_mem[ 7900] = 0;
disk_mem[ 7901] = 0;
disk_mem[ 7902] = 0;
disk_mem[ 7903] = 0;
disk_mem[ 7904] = 0;
disk_mem[ 7905] = 0;
disk_mem[ 7906] = 0;
disk_mem[ 7907] = 0;
disk_mem[ 7908] = 0;
disk_mem[ 7909] = 0;
disk_mem[ 7910] = 0;
disk_mem[ 7911] = 0;
disk_mem[ 7912] = 0;
disk_mem[ 7913] = 0;
disk_mem[ 7914] = 0;
disk_mem[ 7915] = 0;
disk_mem[ 7916] = 0;
disk_mem[ 7917] = 0;
disk_mem[ 7918] = 0;
disk_mem[ 7919] = 0;
disk_mem[ 7920] = 0;
disk_mem[ 7921] = 0;
disk_mem[ 7922] = 0;
disk_mem[ 7923] = 0;
disk_mem[ 7924] = 0;
disk_mem[ 7925] = 0;
disk_mem[ 7926] = 0;
disk_mem[ 7927] = 0;
disk_mem[ 7928] = 0;
disk_mem[ 7929] = 0;
disk_mem[ 7930] = 0;
disk_mem[ 7931] = 0;
disk_mem[ 7932] = 0;
disk_mem[ 7933] = 0;
disk_mem[ 7934] = 0;
disk_mem[ 7935] = 0;
disk_mem[ 7936] = 0;
disk_mem[ 7937] = 0;
disk_mem[ 7938] = 0;
disk_mem[ 7939] = 0;
disk_mem[ 7940] = 0;
disk_mem[ 7941] = 0;
disk_mem[ 7942] = 0;
disk_mem[ 7943] = 0;
disk_mem[ 7944] = 0;
disk_mem[ 7945] = 0;
disk_mem[ 7946] = 0;
disk_mem[ 7947] = 0;
disk_mem[ 7948] = 0;
disk_mem[ 7949] = 0;
disk_mem[ 7950] = 0;
disk_mem[ 7951] = 0;
disk_mem[ 7952] = 0;
disk_mem[ 7953] = 0;
disk_mem[ 7954] = 0;
disk_mem[ 7955] = 0;
disk_mem[ 7956] = 0;
disk_mem[ 7957] = 0;
disk_mem[ 7958] = 0;
disk_mem[ 7959] = 0;
disk_mem[ 7960] = 0;
disk_mem[ 7961] = 0;
disk_mem[ 7962] = 0;
disk_mem[ 7963] = 0;
disk_mem[ 7964] = 0;
disk_mem[ 7965] = 0;
disk_mem[ 7966] = 0;
disk_mem[ 7967] = 0;
disk_mem[ 7968] = 0;
disk_mem[ 7969] = 0;
disk_mem[ 7970] = 0;
disk_mem[ 7971] = 0;
disk_mem[ 7972] = 0;
disk_mem[ 7973] = 0;
disk_mem[ 7974] = 0;
disk_mem[ 7975] = 0;
disk_mem[ 7976] = 0;
disk_mem[ 7977] = 0;
disk_mem[ 7978] = 0;
disk_mem[ 7979] = 0;
disk_mem[ 7980] = 0;
disk_mem[ 7981] = 0;
disk_mem[ 7982] = 0;
disk_mem[ 7983] = 0;
disk_mem[ 7984] = 0;
disk_mem[ 7985] = 0;
disk_mem[ 7986] = 0;
disk_mem[ 7987] = 0;
disk_mem[ 7988] = 0;
disk_mem[ 7989] = 0;
disk_mem[ 7990] = 0;
disk_mem[ 7991] = 0;
disk_mem[ 7992] = 0;
disk_mem[ 7993] = 0;
disk_mem[ 7994] = 0;
disk_mem[ 7995] = 0;
disk_mem[ 7996] = 0;
disk_mem[ 7997] = 0;
disk_mem[ 7998] = 0;
disk_mem[ 7999] = 0;
disk_mem[ 8000] = 0;
disk_mem[ 8001] = 0;
disk_mem[ 8002] = 0;
disk_mem[ 8003] = 0;
disk_mem[ 8004] = 0;
disk_mem[ 8005] = 0;
disk_mem[ 8006] = 0;
disk_mem[ 8007] = 0;
disk_mem[ 8008] = 0;
disk_mem[ 8009] = 0;
disk_mem[ 8010] = 0;
disk_mem[ 8011] = 0;
disk_mem[ 8012] = 0;
disk_mem[ 8013] = 0;
disk_mem[ 8014] = 0;
disk_mem[ 8015] = 0;
disk_mem[ 8016] = 0;
disk_mem[ 8017] = 0;
disk_mem[ 8018] = 0;
disk_mem[ 8019] = 0;
disk_mem[ 8020] = 0;
disk_mem[ 8021] = 0;
disk_mem[ 8022] = 0;
disk_mem[ 8023] = 0;
disk_mem[ 8024] = 0;
disk_mem[ 8025] = 0;
disk_mem[ 8026] = 0;
disk_mem[ 8027] = 0;
disk_mem[ 8028] = 0;
disk_mem[ 8029] = 0;
disk_mem[ 8030] = 0;
disk_mem[ 8031] = 0;
disk_mem[ 8032] = 0;
disk_mem[ 8033] = 0;
disk_mem[ 8034] = 0;
disk_mem[ 8035] = 0;
disk_mem[ 8036] = 0;
disk_mem[ 8037] = 0;
disk_mem[ 8038] = 0;
disk_mem[ 8039] = 0;
disk_mem[ 8040] = 0;
disk_mem[ 8041] = 0;
disk_mem[ 8042] = 0;
disk_mem[ 8043] = 0;
disk_mem[ 8044] = 0;
disk_mem[ 8045] = 0;
disk_mem[ 8046] = 0;
disk_mem[ 8047] = 0;
disk_mem[ 8048] = 0;
disk_mem[ 8049] = 0;
disk_mem[ 8050] = 0;
disk_mem[ 8051] = 0;
disk_mem[ 8052] = 0;
disk_mem[ 8053] = 0;
disk_mem[ 8054] = 0;
disk_mem[ 8055] = 0;
disk_mem[ 8056] = 0;
disk_mem[ 8057] = 0;
disk_mem[ 8058] = 0;
disk_mem[ 8059] = 0;
disk_mem[ 8060] = 0;
disk_mem[ 8061] = 0;
disk_mem[ 8062] = 0;
disk_mem[ 8063] = 0;
disk_mem[ 8064] = 0;
disk_mem[ 8065] = 0;
disk_mem[ 8066] = 0;
disk_mem[ 8067] = 0;
disk_mem[ 8068] = 0;
disk_mem[ 8069] = 0;
disk_mem[ 8070] = 0;
disk_mem[ 8071] = 0;
disk_mem[ 8072] = 0;
disk_mem[ 8073] = 0;
disk_mem[ 8074] = 0;
disk_mem[ 8075] = 0;
disk_mem[ 8076] = 0;
disk_mem[ 8077] = 0;
disk_mem[ 8078] = 0;
disk_mem[ 8079] = 0;
disk_mem[ 8080] = 0;
disk_mem[ 8081] = 0;
disk_mem[ 8082] = 0;
disk_mem[ 8083] = 0;
disk_mem[ 8084] = 0;
disk_mem[ 8085] = 0;
disk_mem[ 8086] = 0;
disk_mem[ 8087] = 0;
disk_mem[ 8088] = 0;
disk_mem[ 8089] = 0;
disk_mem[ 8090] = 0;
disk_mem[ 8091] = 0;
disk_mem[ 8092] = 0;
disk_mem[ 8093] = 0;
disk_mem[ 8094] = 0;
disk_mem[ 8095] = 0;
disk_mem[ 8096] = 0;
disk_mem[ 8097] = 0;
disk_mem[ 8098] = 0;
disk_mem[ 8099] = 0;
disk_mem[ 8100] = 0;
disk_mem[ 8101] = 0;
disk_mem[ 8102] = 0;
disk_mem[ 8103] = 0;
disk_mem[ 8104] = 0;
disk_mem[ 8105] = 0;
disk_mem[ 8106] = 0;
disk_mem[ 8107] = 0;
disk_mem[ 8108] = 0;
disk_mem[ 8109] = 0;
disk_mem[ 8110] = 0;
disk_mem[ 8111] = 0;
disk_mem[ 8112] = 0;
disk_mem[ 8113] = 0;
disk_mem[ 8114] = 0;
disk_mem[ 8115] = 0;
disk_mem[ 8116] = 0;
disk_mem[ 8117] = 0;
disk_mem[ 8118] = 0;
disk_mem[ 8119] = 0;
disk_mem[ 8120] = 0;
disk_mem[ 8121] = 0;
disk_mem[ 8122] = 0;
disk_mem[ 8123] = 0;
disk_mem[ 8124] = 0;
disk_mem[ 8125] = 0;
disk_mem[ 8126] = 0;
disk_mem[ 8127] = 0;
disk_mem[ 8128] = 0;
disk_mem[ 8129] = 0;
disk_mem[ 8130] = 0;
disk_mem[ 8131] = 0;
disk_mem[ 8132] = 0;
disk_mem[ 8133] = 0;
disk_mem[ 8134] = 0;
disk_mem[ 8135] = 0;
disk_mem[ 8136] = 0;
disk_mem[ 8137] = 0;
disk_mem[ 8138] = 0;
disk_mem[ 8139] = 0;
disk_mem[ 8140] = 0;
disk_mem[ 8141] = 0;
disk_mem[ 8142] = 0;
disk_mem[ 8143] = 0;
disk_mem[ 8144] = 0;
disk_mem[ 8145] = 0;
disk_mem[ 8146] = 0;
disk_mem[ 8147] = 0;
disk_mem[ 8148] = 0;
disk_mem[ 8149] = 0;
disk_mem[ 8150] = 0;
disk_mem[ 8151] = 0;
disk_mem[ 8152] = 0;
disk_mem[ 8153] = 0;
disk_mem[ 8154] = 0;
disk_mem[ 8155] = 0;
disk_mem[ 8156] = 0;
disk_mem[ 8157] = 0;
disk_mem[ 8158] = 0;
disk_mem[ 8159] = 0;
disk_mem[ 8160] = 0;
disk_mem[ 8161] = 0;
disk_mem[ 8162] = 0;
disk_mem[ 8163] = 0;
disk_mem[ 8164] = 0;
disk_mem[ 8165] = 0;
disk_mem[ 8166] = 0;
disk_mem[ 8167] = 0;
disk_mem[ 8168] = 0;
disk_mem[ 8169] = 0;
disk_mem[ 8170] = 0;
disk_mem[ 8171] = 0;
disk_mem[ 8172] = 0;
disk_mem[ 8173] = 0;
disk_mem[ 8174] = 0;
disk_mem[ 8175] = 0;
disk_mem[ 8176] = 0;
disk_mem[ 8177] = 0;
disk_mem[ 8178] = 0;
disk_mem[ 8179] = 0;
disk_mem[ 8180] = 0;
disk_mem[ 8181] = 0;
disk_mem[ 8182] = 0;
disk_mem[ 8183] = 0;
disk_mem[ 8184] = 0;
disk_mem[ 8185] = 0;
disk_mem[ 8186] = 0;
disk_mem[ 8187] = 0;
disk_mem[ 8188] = 0;
disk_mem[ 8189] = 0;
disk_mem[ 8190] = 0;
disk_mem[ 8191] = 0;
disk_mem[ 8192] = 0;
disk_mem[ 8193] = 0;
disk_mem[ 8194] = 0;
disk_mem[ 8195] = 0;
disk_mem[ 8196] = 0;
disk_mem[ 8197] = 0;
disk_mem[ 8198] = 0;
disk_mem[ 8199] = 0;
disk_mem[ 8200] = 0;
disk_mem[ 8201] = 0;
disk_mem[ 8202] = 0;
disk_mem[ 8203] = 0;
disk_mem[ 8204] = 0;
disk_mem[ 8205] = 0;
disk_mem[ 8206] = 0;
disk_mem[ 8207] = 0;
disk_mem[ 8208] = 0;
disk_mem[ 8209] = 0;
disk_mem[ 8210] = 0;
disk_mem[ 8211] = 0;
disk_mem[ 8212] = 0;
disk_mem[ 8213] = 0;
disk_mem[ 8214] = 0;
disk_mem[ 8215] = 0;
disk_mem[ 8216] = 0;
disk_mem[ 8217] = 0;
disk_mem[ 8218] = 0;
disk_mem[ 8219] = 0;
disk_mem[ 8220] = 0;
disk_mem[ 8221] = 0;
disk_mem[ 8222] = 0;
disk_mem[ 8223] = 0;
disk_mem[ 8224] = 0;
disk_mem[ 8225] = 0;
disk_mem[ 8226] = 0;
disk_mem[ 8227] = 0;
disk_mem[ 8228] = 0;
disk_mem[ 8229] = 0;
disk_mem[ 8230] = 0;
disk_mem[ 8231] = 0;
disk_mem[ 8232] = 0;
disk_mem[ 8233] = 0;
disk_mem[ 8234] = 0;
disk_mem[ 8235] = 0;
disk_mem[ 8236] = 0;
disk_mem[ 8237] = 0;
disk_mem[ 8238] = 0;
disk_mem[ 8239] = 0;
disk_mem[ 8240] = 0;
disk_mem[ 8241] = 0;
disk_mem[ 8242] = 0;
disk_mem[ 8243] = 0;
disk_mem[ 8244] = 0;
disk_mem[ 8245] = 0;
disk_mem[ 8246] = 0;
disk_mem[ 8247] = 0;
disk_mem[ 8248] = 0;
disk_mem[ 8249] = 0;
disk_mem[ 8250] = 0;
disk_mem[ 8251] = 0;
disk_mem[ 8252] = 0;
disk_mem[ 8253] = 0;
disk_mem[ 8254] = 0;
disk_mem[ 8255] = 0;
disk_mem[ 8256] = 0;
disk_mem[ 8257] = 0;
disk_mem[ 8258] = 0;
disk_mem[ 8259] = 0;
disk_mem[ 8260] = 0;
disk_mem[ 8261] = 0;
disk_mem[ 8262] = 0;
disk_mem[ 8263] = 0;
disk_mem[ 8264] = 0;
disk_mem[ 8265] = 0;
disk_mem[ 8266] = 0;
disk_mem[ 8267] = 0;
disk_mem[ 8268] = 0;
disk_mem[ 8269] = 0;
disk_mem[ 8270] = 0;
disk_mem[ 8271] = 0;
disk_mem[ 8272] = 0;
disk_mem[ 8273] = 0;
disk_mem[ 8274] = 0;
disk_mem[ 8275] = 0;
disk_mem[ 8276] = 0;
disk_mem[ 8277] = 0;
disk_mem[ 8278] = 0;
disk_mem[ 8279] = 0;
disk_mem[ 8280] = 0;
disk_mem[ 8281] = 0;
disk_mem[ 8282] = 0;
disk_mem[ 8283] = 0;
disk_mem[ 8284] = 0;
disk_mem[ 8285] = 0;
disk_mem[ 8286] = 0;
disk_mem[ 8287] = 0;
disk_mem[ 8288] = 0;
disk_mem[ 8289] = 0;
disk_mem[ 8290] = 0;
disk_mem[ 8291] = 0;
disk_mem[ 8292] = 0;
disk_mem[ 8293] = 0;
disk_mem[ 8294] = 0;
disk_mem[ 8295] = 0;
disk_mem[ 8296] = 0;
disk_mem[ 8297] = 0;
disk_mem[ 8298] = 0;
disk_mem[ 8299] = 0;
disk_mem[ 8300] = 0;
disk_mem[ 8301] = 0;
disk_mem[ 8302] = 0;
disk_mem[ 8303] = 0;
disk_mem[ 8304] = 0;
disk_mem[ 8305] = 0;
disk_mem[ 8306] = 0;
disk_mem[ 8307] = 0;
disk_mem[ 8308] = 0;
disk_mem[ 8309] = 0;
disk_mem[ 8310] = 0;
disk_mem[ 8311] = 0;
disk_mem[ 8312] = 0;
disk_mem[ 8313] = 0;
disk_mem[ 8314] = 0;
disk_mem[ 8315] = 0;
disk_mem[ 8316] = 0;
disk_mem[ 8317] = 0;
disk_mem[ 8318] = 0;
disk_mem[ 8319] = 0;
disk_mem[ 8320] = 0;
disk_mem[ 8321] = 0;
disk_mem[ 8322] = 0;
disk_mem[ 8323] = 0;
disk_mem[ 8324] = 0;
disk_mem[ 8325] = 0;
disk_mem[ 8326] = 0;
disk_mem[ 8327] = 0;
disk_mem[ 8328] = 0;
disk_mem[ 8329] = 0;
disk_mem[ 8330] = 0;
disk_mem[ 8331] = 0;
disk_mem[ 8332] = 0;
disk_mem[ 8333] = 0;
disk_mem[ 8334] = 0;
disk_mem[ 8335] = 0;
disk_mem[ 8336] = 0;
disk_mem[ 8337] = 0;
disk_mem[ 8338] = 0;
disk_mem[ 8339] = 0;
disk_mem[ 8340] = 0;
disk_mem[ 8341] = 0;
disk_mem[ 8342] = 0;
disk_mem[ 8343] = 0;
disk_mem[ 8344] = 0;
disk_mem[ 8345] = 0;
disk_mem[ 8346] = 0;
disk_mem[ 8347] = 0;
disk_mem[ 8348] = 0;
disk_mem[ 8349] = 0;
disk_mem[ 8350] = 0;
disk_mem[ 8351] = 0;
disk_mem[ 8352] = 0;
disk_mem[ 8353] = 0;
disk_mem[ 8354] = 0;
disk_mem[ 8355] = 0;
disk_mem[ 8356] = 0;
disk_mem[ 8357] = 0;
disk_mem[ 8358] = 0;
disk_mem[ 8359] = 0;
disk_mem[ 8360] = 0;
disk_mem[ 8361] = 0;
disk_mem[ 8362] = 0;
disk_mem[ 8363] = 0;
disk_mem[ 8364] = 0;
disk_mem[ 8365] = 0;
disk_mem[ 8366] = 0;
disk_mem[ 8367] = 0;
disk_mem[ 8368] = 0;
disk_mem[ 8369] = 0;
disk_mem[ 8370] = 0;
disk_mem[ 8371] = 0;
disk_mem[ 8372] = 0;
disk_mem[ 8373] = 0;
disk_mem[ 8374] = 0;
disk_mem[ 8375] = 0;
disk_mem[ 8376] = 0;
disk_mem[ 8377] = 0;
disk_mem[ 8378] = 0;
disk_mem[ 8379] = 0;
disk_mem[ 8380] = 0;
disk_mem[ 8381] = 0;
disk_mem[ 8382] = 0;
disk_mem[ 8383] = 0;
disk_mem[ 8384] = 0;
disk_mem[ 8385] = 0;
disk_mem[ 8386] = 0;
disk_mem[ 8387] = 0;
disk_mem[ 8388] = 0;
disk_mem[ 8389] = 0;
disk_mem[ 8390] = 0;
disk_mem[ 8391] = 0;
disk_mem[ 8392] = 0;
disk_mem[ 8393] = 0;
disk_mem[ 8394] = 0;
disk_mem[ 8395] = 0;
disk_mem[ 8396] = 0;
disk_mem[ 8397] = 0;
disk_mem[ 8398] = 0;
disk_mem[ 8399] = 0;
disk_mem[ 8400] = 0;
disk_mem[ 8401] = 0;
disk_mem[ 8402] = 0;
disk_mem[ 8403] = 0;
disk_mem[ 8404] = 0;
disk_mem[ 8405] = 0;
disk_mem[ 8406] = 0;
disk_mem[ 8407] = 0;
disk_mem[ 8408] = 0;
disk_mem[ 8409] = 0;
disk_mem[ 8410] = 0;
disk_mem[ 8411] = 0;
disk_mem[ 8412] = 0;
disk_mem[ 8413] = 0;
disk_mem[ 8414] = 0;
disk_mem[ 8415] = 0;
disk_mem[ 8416] = 0;
disk_mem[ 8417] = 0;
disk_mem[ 8418] = 0;
disk_mem[ 8419] = 0;
disk_mem[ 8420] = 0;
disk_mem[ 8421] = 0;
disk_mem[ 8422] = 0;
disk_mem[ 8423] = 0;
disk_mem[ 8424] = 0;
disk_mem[ 8425] = 0;
disk_mem[ 8426] = 0;
disk_mem[ 8427] = 0;
disk_mem[ 8428] = 0;
disk_mem[ 8429] = 0;
disk_mem[ 8430] = 0;
disk_mem[ 8431] = 0;
disk_mem[ 8432] = 0;
disk_mem[ 8433] = 0;
disk_mem[ 8434] = 0;
disk_mem[ 8435] = 0;
disk_mem[ 8436] = 0;
disk_mem[ 8437] = 0;
disk_mem[ 8438] = 0;
disk_mem[ 8439] = 0;
disk_mem[ 8440] = 0;
disk_mem[ 8441] = 0;
disk_mem[ 8442] = 0;
disk_mem[ 8443] = 0;
disk_mem[ 8444] = 0;
disk_mem[ 8445] = 0;
disk_mem[ 8446] = 0;
disk_mem[ 8447] = 0;
disk_mem[ 8448] = 0;
disk_mem[ 8449] = 0;
disk_mem[ 8450] = 0;
disk_mem[ 8451] = 0;
disk_mem[ 8452] = 0;
disk_mem[ 8453] = 0;
disk_mem[ 8454] = 0;
disk_mem[ 8455] = 0;
disk_mem[ 8456] = 0;
disk_mem[ 8457] = 0;
disk_mem[ 8458] = 0;
disk_mem[ 8459] = 0;
disk_mem[ 8460] = 0;
disk_mem[ 8461] = 0;
disk_mem[ 8462] = 0;
disk_mem[ 8463] = 0;
disk_mem[ 8464] = 0;
disk_mem[ 8465] = 0;
disk_mem[ 8466] = 0;
disk_mem[ 8467] = 0;
disk_mem[ 8468] = 0;
disk_mem[ 8469] = 0;
disk_mem[ 8470] = 0;
disk_mem[ 8471] = 0;
disk_mem[ 8472] = 0;
disk_mem[ 8473] = 0;
disk_mem[ 8474] = 0;
disk_mem[ 8475] = 0;
disk_mem[ 8476] = 0;
disk_mem[ 8477] = 0;
disk_mem[ 8478] = 0;
disk_mem[ 8479] = 0;
disk_mem[ 8480] = 0;
disk_mem[ 8481] = 0;
disk_mem[ 8482] = 0;
disk_mem[ 8483] = 0;
disk_mem[ 8484] = 0;
disk_mem[ 8485] = 0;
disk_mem[ 8486] = 0;
disk_mem[ 8487] = 0;
disk_mem[ 8488] = 0;
disk_mem[ 8489] = 0;
disk_mem[ 8490] = 0;
disk_mem[ 8491] = 0;
disk_mem[ 8492] = 0;
disk_mem[ 8493] = 0;
disk_mem[ 8494] = 0;
disk_mem[ 8495] = 0;
disk_mem[ 8496] = 0;
disk_mem[ 8497] = 0;
disk_mem[ 8498] = 0;
disk_mem[ 8499] = 0;
disk_mem[ 8500] = 0;
disk_mem[ 8501] = 0;
disk_mem[ 8502] = 0;
disk_mem[ 8503] = 0;
disk_mem[ 8504] = 0;
disk_mem[ 8505] = 0;
disk_mem[ 8506] = 0;
disk_mem[ 8507] = 0;
disk_mem[ 8508] = 0;
disk_mem[ 8509] = 0;
disk_mem[ 8510] = 0;
disk_mem[ 8511] = 0;
disk_mem[ 8512] = 0;
disk_mem[ 8513] = 0;
disk_mem[ 8514] = 0;
disk_mem[ 8515] = 0;
disk_mem[ 8516] = 0;
disk_mem[ 8517] = 0;
disk_mem[ 8518] = 0;
disk_mem[ 8519] = 0;
disk_mem[ 8520] = 0;
disk_mem[ 8521] = 0;
disk_mem[ 8522] = 0;
disk_mem[ 8523] = 0;
disk_mem[ 8524] = 0;
disk_mem[ 8525] = 0;
disk_mem[ 8526] = 0;
disk_mem[ 8527] = 0;
disk_mem[ 8528] = 0;
disk_mem[ 8529] = 0;
disk_mem[ 8530] = 0;
disk_mem[ 8531] = 0;
disk_mem[ 8532] = 0;
disk_mem[ 8533] = 0;
disk_mem[ 8534] = 0;
disk_mem[ 8535] = 0;
disk_mem[ 8536] = 0;
disk_mem[ 8537] = 0;
disk_mem[ 8538] = 0;
disk_mem[ 8539] = 0;
disk_mem[ 8540] = 0;
disk_mem[ 8541] = 0;
disk_mem[ 8542] = 0;
disk_mem[ 8543] = 0;
disk_mem[ 8544] = 0;
disk_mem[ 8545] = 0;
disk_mem[ 8546] = 0;
disk_mem[ 8547] = 0;
disk_mem[ 8548] = 0;
disk_mem[ 8549] = 0;
disk_mem[ 8550] = 0;
disk_mem[ 8551] = 0;
disk_mem[ 8552] = 0;
disk_mem[ 8553] = 0;
disk_mem[ 8554] = 0;
disk_mem[ 8555] = 0;
disk_mem[ 8556] = 0;
disk_mem[ 8557] = 0;
disk_mem[ 8558] = 0;
disk_mem[ 8559] = 0;
disk_mem[ 8560] = 0;
disk_mem[ 8561] = 0;
disk_mem[ 8562] = 0;
disk_mem[ 8563] = 0;
disk_mem[ 8564] = 0;
disk_mem[ 8565] = 0;
disk_mem[ 8566] = 0;
disk_mem[ 8567] = 0;
disk_mem[ 8568] = 0;
disk_mem[ 8569] = 0;
disk_mem[ 8570] = 0;
disk_mem[ 8571] = 0;
disk_mem[ 8572] = 0;
disk_mem[ 8573] = 0;
disk_mem[ 8574] = 0;
disk_mem[ 8575] = 0;
disk_mem[ 8576] = 0;
disk_mem[ 8577] = 0;
disk_mem[ 8578] = 0;
disk_mem[ 8579] = 0;
disk_mem[ 8580] = 0;
disk_mem[ 8581] = 0;
disk_mem[ 8582] = 0;
disk_mem[ 8583] = 0;
disk_mem[ 8584] = 0;
disk_mem[ 8585] = 0;
disk_mem[ 8586] = 0;
disk_mem[ 8587] = 0;
disk_mem[ 8588] = 0;
disk_mem[ 8589] = 0;
disk_mem[ 8590] = 0;
disk_mem[ 8591] = 0;
disk_mem[ 8592] = 0;
disk_mem[ 8593] = 0;
disk_mem[ 8594] = 0;
disk_mem[ 8595] = 0;
disk_mem[ 8596] = 0;
disk_mem[ 8597] = 0;
disk_mem[ 8598] = 0;
disk_mem[ 8599] = 0;
disk_mem[ 8600] = 0;
disk_mem[ 8601] = 0;
disk_mem[ 8602] = 0;
disk_mem[ 8603] = 0;
disk_mem[ 8604] = 0;
disk_mem[ 8605] = 0;
disk_mem[ 8606] = 0;
disk_mem[ 8607] = 0;
disk_mem[ 8608] = 0;
disk_mem[ 8609] = 0;
disk_mem[ 8610] = 0;
disk_mem[ 8611] = 0;
disk_mem[ 8612] = 0;
disk_mem[ 8613] = 0;
disk_mem[ 8614] = 0;
disk_mem[ 8615] = 0;
disk_mem[ 8616] = 0;
disk_mem[ 8617] = 0;
disk_mem[ 8618] = 0;
disk_mem[ 8619] = 0;
disk_mem[ 8620] = 0;
disk_mem[ 8621] = 0;
disk_mem[ 8622] = 0;
disk_mem[ 8623] = 0;
disk_mem[ 8624] = 0;
disk_mem[ 8625] = 0;
disk_mem[ 8626] = 0;
disk_mem[ 8627] = 0;
disk_mem[ 8628] = 0;
disk_mem[ 8629] = 0;
disk_mem[ 8630] = 0;
disk_mem[ 8631] = 0;
disk_mem[ 8632] = 0;
disk_mem[ 8633] = 0;
disk_mem[ 8634] = 0;
disk_mem[ 8635] = 0;
disk_mem[ 8636] = 0;
disk_mem[ 8637] = 0;
disk_mem[ 8638] = 0;
disk_mem[ 8639] = 0;
disk_mem[ 8640] = 0;
disk_mem[ 8641] = 0;
disk_mem[ 8642] = 0;
disk_mem[ 8643] = 0;
disk_mem[ 8644] = 0;
disk_mem[ 8645] = 0;
disk_mem[ 8646] = 0;
disk_mem[ 8647] = 0;
disk_mem[ 8648] = 0;
disk_mem[ 8649] = 0;
disk_mem[ 8650] = 0;
disk_mem[ 8651] = 0;
disk_mem[ 8652] = 0;
disk_mem[ 8653] = 0;
disk_mem[ 8654] = 0;
disk_mem[ 8655] = 0;
disk_mem[ 8656] = 0;
disk_mem[ 8657] = 0;
disk_mem[ 8658] = 0;
disk_mem[ 8659] = 0;
disk_mem[ 8660] = 0;
disk_mem[ 8661] = 0;
disk_mem[ 8662] = 0;
disk_mem[ 8663] = 0;
disk_mem[ 8664] = 0;
disk_mem[ 8665] = 0;
disk_mem[ 8666] = 0;
disk_mem[ 8667] = 0;
disk_mem[ 8668] = 0;
disk_mem[ 8669] = 0;
disk_mem[ 8670] = 0;
disk_mem[ 8671] = 0;
disk_mem[ 8672] = 0;
disk_mem[ 8673] = 0;
disk_mem[ 8674] = 0;
disk_mem[ 8675] = 0;
disk_mem[ 8676] = 0;
disk_mem[ 8677] = 0;
disk_mem[ 8678] = 0;
disk_mem[ 8679] = 0;
disk_mem[ 8680] = 0;
disk_mem[ 8681] = 0;
disk_mem[ 8682] = 0;
disk_mem[ 8683] = 0;
disk_mem[ 8684] = 0;
disk_mem[ 8685] = 0;
disk_mem[ 8686] = 0;
disk_mem[ 8687] = 0;
disk_mem[ 8688] = 0;
disk_mem[ 8689] = 0;
disk_mem[ 8690] = 0;
disk_mem[ 8691] = 0;
disk_mem[ 8692] = 0;
disk_mem[ 8693] = 0;
disk_mem[ 8694] = 0;
disk_mem[ 8695] = 0;
disk_mem[ 8696] = 0;
disk_mem[ 8697] = 0;
disk_mem[ 8698] = 0;
disk_mem[ 8699] = 0;
disk_mem[ 8700] = 0;
disk_mem[ 8701] = 0;
disk_mem[ 8702] = 0;
disk_mem[ 8703] = 0;
disk_mem[ 8704] = 0;
disk_mem[ 8705] = 0;
disk_mem[ 8706] = 0;
disk_mem[ 8707] = 0;
disk_mem[ 8708] = 0;
disk_mem[ 8709] = 0;
disk_mem[ 8710] = 0;
disk_mem[ 8711] = 0;
disk_mem[ 8712] = 0;
disk_mem[ 8713] = 0;
disk_mem[ 8714] = 0;
disk_mem[ 8715] = 0;
disk_mem[ 8716] = 0;
disk_mem[ 8717] = 0;
disk_mem[ 8718] = 0;
disk_mem[ 8719] = 0;
disk_mem[ 8720] = 0;
disk_mem[ 8721] = 0;
disk_mem[ 8722] = 0;
disk_mem[ 8723] = 0;
disk_mem[ 8724] = 0;
disk_mem[ 8725] = 0;
disk_mem[ 8726] = 0;
disk_mem[ 8727] = 0;
disk_mem[ 8728] = 0;
disk_mem[ 8729] = 0;
disk_mem[ 8730] = 0;
disk_mem[ 8731] = 0;
disk_mem[ 8732] = 0;
disk_mem[ 8733] = 0;
disk_mem[ 8734] = 0;
disk_mem[ 8735] = 0;
disk_mem[ 8736] = 0;
disk_mem[ 8737] = 0;
disk_mem[ 8738] = 0;
disk_mem[ 8739] = 0;
disk_mem[ 8740] = 0;
disk_mem[ 8741] = 0;
disk_mem[ 8742] = 0;
disk_mem[ 8743] = 0;
disk_mem[ 8744] = 0;
disk_mem[ 8745] = 0;
disk_mem[ 8746] = 0;
disk_mem[ 8747] = 0;
disk_mem[ 8748] = 0;
disk_mem[ 8749] = 0;
disk_mem[ 8750] = 0;
disk_mem[ 8751] = 0;
disk_mem[ 8752] = 0;
disk_mem[ 8753] = 0;
disk_mem[ 8754] = 0;
disk_mem[ 8755] = 0;
disk_mem[ 8756] = 0;
disk_mem[ 8757] = 0;
disk_mem[ 8758] = 0;
disk_mem[ 8759] = 0;
disk_mem[ 8760] = 0;
disk_mem[ 8761] = 0;
disk_mem[ 8762] = 0;
disk_mem[ 8763] = 0;
disk_mem[ 8764] = 0;
disk_mem[ 8765] = 0;
disk_mem[ 8766] = 0;
disk_mem[ 8767] = 0;
disk_mem[ 8768] = 0;
disk_mem[ 8769] = 0;
disk_mem[ 8770] = 0;
disk_mem[ 8771] = 0;
disk_mem[ 8772] = 0;
disk_mem[ 8773] = 0;
disk_mem[ 8774] = 0;
disk_mem[ 8775] = 0;
disk_mem[ 8776] = 0;
disk_mem[ 8777] = 0;
disk_mem[ 8778] = 0;
disk_mem[ 8779] = 0;
disk_mem[ 8780] = 0;
disk_mem[ 8781] = 0;
disk_mem[ 8782] = 0;
disk_mem[ 8783] = 0;
disk_mem[ 8784] = 0;
disk_mem[ 8785] = 0;
disk_mem[ 8786] = 0;
disk_mem[ 8787] = 0;
disk_mem[ 8788] = 0;
disk_mem[ 8789] = 0;
disk_mem[ 8790] = 0;
disk_mem[ 8791] = 0;
disk_mem[ 8792] = 0;
disk_mem[ 8793] = 0;
disk_mem[ 8794] = 0;
disk_mem[ 8795] = 0;
disk_mem[ 8796] = 0;
disk_mem[ 8797] = 0;
disk_mem[ 8798] = 0;
disk_mem[ 8799] = 0;
disk_mem[ 8800] = 0;
disk_mem[ 8801] = 0;
disk_mem[ 8802] = 0;
disk_mem[ 8803] = 0;
disk_mem[ 8804] = 0;
disk_mem[ 8805] = 0;
disk_mem[ 8806] = 0;
disk_mem[ 8807] = 0;
disk_mem[ 8808] = 0;
disk_mem[ 8809] = 0;
disk_mem[ 8810] = 0;
disk_mem[ 8811] = 0;
disk_mem[ 8812] = 0;
disk_mem[ 8813] = 0;
disk_mem[ 8814] = 0;
disk_mem[ 8815] = 0;
disk_mem[ 8816] = 0;
disk_mem[ 8817] = 0;
disk_mem[ 8818] = 0;
disk_mem[ 8819] = 0;
disk_mem[ 8820] = 0;
disk_mem[ 8821] = 0;
disk_mem[ 8822] = 0;
disk_mem[ 8823] = 0;
disk_mem[ 8824] = 0;
disk_mem[ 8825] = 0;
disk_mem[ 8826] = 0;
disk_mem[ 8827] = 0;
disk_mem[ 8828] = 0;
disk_mem[ 8829] = 0;
disk_mem[ 8830] = 0;
disk_mem[ 8831] = 0;
disk_mem[ 8832] = 0;
disk_mem[ 8833] = 0;
disk_mem[ 8834] = 0;
disk_mem[ 8835] = 0;
disk_mem[ 8836] = 0;
disk_mem[ 8837] = 0;
disk_mem[ 8838] = 0;
disk_mem[ 8839] = 0;
disk_mem[ 8840] = 0;
disk_mem[ 8841] = 0;
disk_mem[ 8842] = 0;
disk_mem[ 8843] = 0;
disk_mem[ 8844] = 0;
disk_mem[ 8845] = 0;
disk_mem[ 8846] = 0;
disk_mem[ 8847] = 0;
disk_mem[ 8848] = 0;
disk_mem[ 8849] = 0;
disk_mem[ 8850] = 0;
disk_mem[ 8851] = 0;
disk_mem[ 8852] = 0;
disk_mem[ 8853] = 0;
disk_mem[ 8854] = 0;
disk_mem[ 8855] = 0;
disk_mem[ 8856] = 0;
disk_mem[ 8857] = 0;
disk_mem[ 8858] = 0;
disk_mem[ 8859] = 0;
disk_mem[ 8860] = 0;
disk_mem[ 8861] = 0;
disk_mem[ 8862] = 0;
disk_mem[ 8863] = 0;
disk_mem[ 8864] = 0;
disk_mem[ 8865] = 0;
disk_mem[ 8866] = 0;
disk_mem[ 8867] = 0;
disk_mem[ 8868] = 0;
disk_mem[ 8869] = 0;
disk_mem[ 8870] = 0;
disk_mem[ 8871] = 0;
disk_mem[ 8872] = 0;
disk_mem[ 8873] = 0;
disk_mem[ 8874] = 0;
disk_mem[ 8875] = 0;
disk_mem[ 8876] = 0;
disk_mem[ 8877] = 0;
disk_mem[ 8878] = 0;
disk_mem[ 8879] = 0;
disk_mem[ 8880] = 0;
disk_mem[ 8881] = 0;
disk_mem[ 8882] = 0;
disk_mem[ 8883] = 0;
disk_mem[ 8884] = 0;
disk_mem[ 8885] = 0;
disk_mem[ 8886] = 0;
disk_mem[ 8887] = 0;
disk_mem[ 8888] = 0;
disk_mem[ 8889] = 0;
disk_mem[ 8890] = 0;
disk_mem[ 8891] = 0;
disk_mem[ 8892] = 0;
disk_mem[ 8893] = 0;
disk_mem[ 8894] = 0;
disk_mem[ 8895] = 0;
disk_mem[ 8896] = 0;
disk_mem[ 8897] = 0;
disk_mem[ 8898] = 0;
disk_mem[ 8899] = 0;
disk_mem[ 8900] = 0;
disk_mem[ 8901] = 0;
disk_mem[ 8902] = 0;
disk_mem[ 8903] = 0;
disk_mem[ 8904] = 0;
disk_mem[ 8905] = 0;
disk_mem[ 8906] = 0;
disk_mem[ 8907] = 0;
disk_mem[ 8908] = 0;
disk_mem[ 8909] = 0;
disk_mem[ 8910] = 0;
disk_mem[ 8911] = 0;
disk_mem[ 8912] = 0;
disk_mem[ 8913] = 0;
disk_mem[ 8914] = 0;
disk_mem[ 8915] = 0;
disk_mem[ 8916] = 0;
disk_mem[ 8917] = 0;
disk_mem[ 8918] = 0;
disk_mem[ 8919] = 0;
disk_mem[ 8920] = 0;
disk_mem[ 8921] = 0;
disk_mem[ 8922] = 0;
disk_mem[ 8923] = 0;
disk_mem[ 8924] = 0;
disk_mem[ 8925] = 0;
disk_mem[ 8926] = 0;
disk_mem[ 8927] = 0;
disk_mem[ 8928] = 0;
disk_mem[ 8929] = 0;
disk_mem[ 8930] = 0;
disk_mem[ 8931] = 0;
disk_mem[ 8932] = 0;
disk_mem[ 8933] = 0;
disk_mem[ 8934] = 0;
disk_mem[ 8935] = 0;
disk_mem[ 8936] = 0;
disk_mem[ 8937] = 0;
disk_mem[ 8938] = 0;
disk_mem[ 8939] = 0;
disk_mem[ 8940] = 0;
disk_mem[ 8941] = 0;
disk_mem[ 8942] = 0;
disk_mem[ 8943] = 0;
disk_mem[ 8944] = 0;
disk_mem[ 8945] = 0;
disk_mem[ 8946] = 0;
disk_mem[ 8947] = 0;
disk_mem[ 8948] = 0;
disk_mem[ 8949] = 0;
disk_mem[ 8950] = 0;
disk_mem[ 8951] = 0;
disk_mem[ 8952] = 0;
disk_mem[ 8953] = 0;
disk_mem[ 8954] = 0;
disk_mem[ 8955] = 0;
disk_mem[ 8956] = 0;
disk_mem[ 8957] = 0;
disk_mem[ 8958] = 0;
disk_mem[ 8959] = 0;
disk_mem[ 8960] = 0;
disk_mem[ 8961] = 0;
disk_mem[ 8962] = 0;
disk_mem[ 8963] = 0;
disk_mem[ 8964] = 0;
disk_mem[ 8965] = 0;
disk_mem[ 8966] = 0;
disk_mem[ 8967] = 0;
disk_mem[ 8968] = 0;
disk_mem[ 8969] = 0;
disk_mem[ 8970] = 0;
disk_mem[ 8971] = 0;
disk_mem[ 8972] = 0;
disk_mem[ 8973] = 0;
disk_mem[ 8974] = 0;
disk_mem[ 8975] = 0;
disk_mem[ 8976] = 0;
disk_mem[ 8977] = 0;
disk_mem[ 8978] = 0;
disk_mem[ 8979] = 0;
disk_mem[ 8980] = 0;
disk_mem[ 8981] = 0;
disk_mem[ 8982] = 0;
disk_mem[ 8983] = 0;
disk_mem[ 8984] = 0;
disk_mem[ 8985] = 0;
disk_mem[ 8986] = 0;
disk_mem[ 8987] = 0;
disk_mem[ 8988] = 0;
disk_mem[ 8989] = 0;
disk_mem[ 8990] = 0;
disk_mem[ 8991] = 0;
disk_mem[ 8992] = 0;
disk_mem[ 8993] = 0;
disk_mem[ 8994] = 0;
disk_mem[ 8995] = 0;
disk_mem[ 8996] = 0;
disk_mem[ 8997] = 0;
disk_mem[ 8998] = 0;
disk_mem[ 8999] = 0;
disk_mem[ 9000] = 0;
disk_mem[ 9001] = 0;
disk_mem[ 9002] = 0;
disk_mem[ 9003] = 0;
disk_mem[ 9004] = 0;
disk_mem[ 9005] = 0;
disk_mem[ 9006] = 0;
disk_mem[ 9007] = 0;
disk_mem[ 9008] = 0;
disk_mem[ 9009] = 0;
disk_mem[ 9010] = 0;
disk_mem[ 9011] = 0;
disk_mem[ 9012] = 0;
disk_mem[ 9013] = 0;
disk_mem[ 9014] = 0;
disk_mem[ 9015] = 0;
disk_mem[ 9016] = 0;
disk_mem[ 9017] = 0;
disk_mem[ 9018] = 0;
disk_mem[ 9019] = 0;
disk_mem[ 9020] = 0;
disk_mem[ 9021] = 0;
disk_mem[ 9022] = 0;
disk_mem[ 9023] = 0;
disk_mem[ 9024] = 0;
disk_mem[ 9025] = 0;
disk_mem[ 9026] = 0;
disk_mem[ 9027] = 0;
disk_mem[ 9028] = 0;
disk_mem[ 9029] = 0;
disk_mem[ 9030] = 0;
disk_mem[ 9031] = 0;
disk_mem[ 9032] = 0;
disk_mem[ 9033] = 0;
disk_mem[ 9034] = 0;
disk_mem[ 9035] = 0;
disk_mem[ 9036] = 0;
disk_mem[ 9037] = 0;
disk_mem[ 9038] = 0;
disk_mem[ 9039] = 0;
disk_mem[ 9040] = 0;
disk_mem[ 9041] = 0;
disk_mem[ 9042] = 0;
disk_mem[ 9043] = 0;
disk_mem[ 9044] = 0;
disk_mem[ 9045] = 0;
disk_mem[ 9046] = 0;
disk_mem[ 9047] = 0;
disk_mem[ 9048] = 0;
disk_mem[ 9049] = 0;
disk_mem[ 9050] = 0;
disk_mem[ 9051] = 0;
disk_mem[ 9052] = 0;
disk_mem[ 9053] = 0;
disk_mem[ 9054] = 0;
disk_mem[ 9055] = 0;
disk_mem[ 9056] = 0;
disk_mem[ 9057] = 0;
disk_mem[ 9058] = 0;
disk_mem[ 9059] = 0;
disk_mem[ 9060] = 0;
disk_mem[ 9061] = 0;
disk_mem[ 9062] = 0;
disk_mem[ 9063] = 0;
disk_mem[ 9064] = 0;
disk_mem[ 9065] = 0;
disk_mem[ 9066] = 0;
disk_mem[ 9067] = 0;
disk_mem[ 9068] = 0;
disk_mem[ 9069] = 0;
disk_mem[ 9070] = 0;
disk_mem[ 9071] = 0;
disk_mem[ 9072] = 0;
disk_mem[ 9073] = 0;
disk_mem[ 9074] = 0;
disk_mem[ 9075] = 0;
disk_mem[ 9076] = 0;
disk_mem[ 9077] = 0;
disk_mem[ 9078] = 0;
disk_mem[ 9079] = 0;
disk_mem[ 9080] = 0;
disk_mem[ 9081] = 0;
disk_mem[ 9082] = 0;
disk_mem[ 9083] = 0;
disk_mem[ 9084] = 0;
disk_mem[ 9085] = 0;
disk_mem[ 9086] = 0;
disk_mem[ 9087] = 0;
disk_mem[ 9088] = 0;
disk_mem[ 9089] = 0;
disk_mem[ 9090] = 0;
disk_mem[ 9091] = 0;
disk_mem[ 9092] = 0;
disk_mem[ 9093] = 0;
disk_mem[ 9094] = 0;
disk_mem[ 9095] = 0;
disk_mem[ 9096] = 0;
disk_mem[ 9097] = 0;
disk_mem[ 9098] = 0;
disk_mem[ 9099] = 0;
disk_mem[ 9100] = 0;
disk_mem[ 9101] = 0;
disk_mem[ 9102] = 0;
disk_mem[ 9103] = 0;
disk_mem[ 9104] = 0;
disk_mem[ 9105] = 0;
disk_mem[ 9106] = 0;
disk_mem[ 9107] = 0;
disk_mem[ 9108] = 0;
disk_mem[ 9109] = 0;
disk_mem[ 9110] = 0;
disk_mem[ 9111] = 0;
disk_mem[ 9112] = 0;
disk_mem[ 9113] = 0;
disk_mem[ 9114] = 0;
disk_mem[ 9115] = 0;
disk_mem[ 9116] = 0;
disk_mem[ 9117] = 0;
disk_mem[ 9118] = 0;
disk_mem[ 9119] = 0;
disk_mem[ 9120] = 0;
disk_mem[ 9121] = 0;
disk_mem[ 9122] = 0;
disk_mem[ 9123] = 0;
disk_mem[ 9124] = 0;
disk_mem[ 9125] = 0;
disk_mem[ 9126] = 0;
disk_mem[ 9127] = 0;
disk_mem[ 9128] = 0;
disk_mem[ 9129] = 0;
disk_mem[ 9130] = 0;
disk_mem[ 9131] = 0;
disk_mem[ 9132] = 0;
disk_mem[ 9133] = 0;
disk_mem[ 9134] = 0;
disk_mem[ 9135] = 0;
disk_mem[ 9136] = 0;
disk_mem[ 9137] = 0;
disk_mem[ 9138] = 0;
disk_mem[ 9139] = 0;
disk_mem[ 9140] = 0;
disk_mem[ 9141] = 0;
disk_mem[ 9142] = 0;
disk_mem[ 9143] = 0;
disk_mem[ 9144] = 0;
disk_mem[ 9145] = 0;
disk_mem[ 9146] = 0;
disk_mem[ 9147] = 0;
disk_mem[ 9148] = 0;
disk_mem[ 9149] = 0;
disk_mem[ 9150] = 0;
disk_mem[ 9151] = 0;
disk_mem[ 9152] = 0;
disk_mem[ 9153] = 0;
disk_mem[ 9154] = 0;
disk_mem[ 9155] = 0;
disk_mem[ 9156] = 0;
disk_mem[ 9157] = 0;
disk_mem[ 9158] = 0;
disk_mem[ 9159] = 0;
disk_mem[ 9160] = 0;
disk_mem[ 9161] = 0;
disk_mem[ 9162] = 0;
disk_mem[ 9163] = 0;
disk_mem[ 9164] = 0;
disk_mem[ 9165] = 0;
disk_mem[ 9166] = 0;
disk_mem[ 9167] = 0;
disk_mem[ 9168] = 0;
disk_mem[ 9169] = 0;
disk_mem[ 9170] = 0;
disk_mem[ 9171] = 0;
disk_mem[ 9172] = 0;
disk_mem[ 9173] = 0;
disk_mem[ 9174] = 0;
disk_mem[ 9175] = 0;
disk_mem[ 9176] = 0;
disk_mem[ 9177] = 0;
disk_mem[ 9178] = 0;
disk_mem[ 9179] = 0;
disk_mem[ 9180] = 0;
disk_mem[ 9181] = 0;
disk_mem[ 9182] = 0;
disk_mem[ 9183] = 0;
disk_mem[ 9184] = 0;
disk_mem[ 9185] = 0;
disk_mem[ 9186] = 0;
disk_mem[ 9187] = 0;
disk_mem[ 9188] = 0;
disk_mem[ 9189] = 0;
disk_mem[ 9190] = 0;
disk_mem[ 9191] = 0;
disk_mem[ 9192] = 0;
disk_mem[ 9193] = 0;
disk_mem[ 9194] = 0;
disk_mem[ 9195] = 0;
disk_mem[ 9196] = 0;
disk_mem[ 9197] = 0;
disk_mem[ 9198] = 0;
disk_mem[ 9199] = 0;
disk_mem[ 9200] = 0;
disk_mem[ 9201] = 0;
disk_mem[ 9202] = 0;
disk_mem[ 9203] = 0;
disk_mem[ 9204] = 0;
disk_mem[ 9205] = 0;
disk_mem[ 9206] = 0;
disk_mem[ 9207] = 0;
disk_mem[ 9208] = 0;
disk_mem[ 9209] = 0;
disk_mem[ 9210] = 0;
disk_mem[ 9211] = 0;
disk_mem[ 9212] = 0;
disk_mem[ 9213] = 0;
disk_mem[ 9214] = 0;
disk_mem[ 9215] = 0;
disk_mem[ 9216] = 0;
disk_mem[ 9217] = 0;
disk_mem[ 9218] = 0;
disk_mem[ 9219] = 0;
disk_mem[ 9220] = 0;
disk_mem[ 9221] = 0;
disk_mem[ 9222] = 0;
disk_mem[ 9223] = 0;
disk_mem[ 9224] = 0;
disk_mem[ 9225] = 0;
disk_mem[ 9226] = 0;
disk_mem[ 9227] = 0;
disk_mem[ 9228] = 0;
disk_mem[ 9229] = 0;
disk_mem[ 9230] = 0;
disk_mem[ 9231] = 0;
disk_mem[ 9232] = 0;
disk_mem[ 9233] = 0;
disk_mem[ 9234] = 0;
disk_mem[ 9235] = 0;
disk_mem[ 9236] = 0;
disk_mem[ 9237] = 0;
disk_mem[ 9238] = 0;
disk_mem[ 9239] = 0;
disk_mem[ 9240] = 0;
disk_mem[ 9241] = 0;
disk_mem[ 9242] = 0;
disk_mem[ 9243] = 0;
disk_mem[ 9244] = 0;
disk_mem[ 9245] = 0;
disk_mem[ 9246] = 0;
disk_mem[ 9247] = 0;
disk_mem[ 9248] = 0;
disk_mem[ 9249] = 0;
disk_mem[ 9250] = 0;
disk_mem[ 9251] = 0;
disk_mem[ 9252] = 0;
disk_mem[ 9253] = 0;
disk_mem[ 9254] = 0;
disk_mem[ 9255] = 0;
disk_mem[ 9256] = 0;
disk_mem[ 9257] = 0;
disk_mem[ 9258] = 0;
disk_mem[ 9259] = 0;
disk_mem[ 9260] = 0;
disk_mem[ 9261] = 0;
disk_mem[ 9262] = 0;
disk_mem[ 9263] = 0;
disk_mem[ 9264] = 0;
disk_mem[ 9265] = 0;
disk_mem[ 9266] = 0;
disk_mem[ 9267] = 0;
disk_mem[ 9268] = 0;
disk_mem[ 9269] = 0;
disk_mem[ 9270] = 0;
disk_mem[ 9271] = 0;
disk_mem[ 9272] = 0;
disk_mem[ 9273] = 0;
disk_mem[ 9274] = 0;
disk_mem[ 9275] = 0;
disk_mem[ 9276] = 0;
disk_mem[ 9277] = 0;
disk_mem[ 9278] = 0;
disk_mem[ 9279] = 0;
disk_mem[ 9280] = 0;
disk_mem[ 9281] = 0;
disk_mem[ 9282] = 0;
disk_mem[ 9283] = 0;
disk_mem[ 9284] = 0;
disk_mem[ 9285] = 0;
disk_mem[ 9286] = 0;
disk_mem[ 9287] = 0;
disk_mem[ 9288] = 0;
disk_mem[ 9289] = 0;
disk_mem[ 9290] = 0;
disk_mem[ 9291] = 0;
disk_mem[ 9292] = 0;
disk_mem[ 9293] = 0;
disk_mem[ 9294] = 0;
disk_mem[ 9295] = 0;
disk_mem[ 9296] = 0;
disk_mem[ 9297] = 0;
disk_mem[ 9298] = 0;
disk_mem[ 9299] = 0;
disk_mem[ 9300] = 0;
disk_mem[ 9301] = 0;
disk_mem[ 9302] = 0;
disk_mem[ 9303] = 0;
disk_mem[ 9304] = 0;
disk_mem[ 9305] = 0;
disk_mem[ 9306] = 0;
disk_mem[ 9307] = 0;
disk_mem[ 9308] = 0;
disk_mem[ 9309] = 0;
disk_mem[ 9310] = 0;
disk_mem[ 9311] = 0;
disk_mem[ 9312] = 0;
disk_mem[ 9313] = 0;
disk_mem[ 9314] = 0;
disk_mem[ 9315] = 0;
disk_mem[ 9316] = 0;
disk_mem[ 9317] = 0;
disk_mem[ 9318] = 0;
disk_mem[ 9319] = 0;
disk_mem[ 9320] = 0;
disk_mem[ 9321] = 0;
disk_mem[ 9322] = 0;
disk_mem[ 9323] = 0;
disk_mem[ 9324] = 0;
disk_mem[ 9325] = 0;
disk_mem[ 9326] = 0;
disk_mem[ 9327] = 0;
disk_mem[ 9328] = 0;
disk_mem[ 9329] = 0;
disk_mem[ 9330] = 0;
disk_mem[ 9331] = 0;
disk_mem[ 9332] = 0;
disk_mem[ 9333] = 0;
disk_mem[ 9334] = 0;
disk_mem[ 9335] = 0;
disk_mem[ 9336] = 0;
disk_mem[ 9337] = 0;
disk_mem[ 9338] = 0;
disk_mem[ 9339] = 0;
disk_mem[ 9340] = 0;
disk_mem[ 9341] = 0;
disk_mem[ 9342] = 0;
disk_mem[ 9343] = 0;
disk_mem[ 9344] = 0;
disk_mem[ 9345] = 0;
disk_mem[ 9346] = 0;
disk_mem[ 9347] = 0;
disk_mem[ 9348] = 0;
disk_mem[ 9349] = 0;
disk_mem[ 9350] = 0;
disk_mem[ 9351] = 0;
disk_mem[ 9352] = 0;
disk_mem[ 9353] = 0;
disk_mem[ 9354] = 0;
disk_mem[ 9355] = 0;
disk_mem[ 9356] = 0;
disk_mem[ 9357] = 0;
disk_mem[ 9358] = 0;
disk_mem[ 9359] = 0;
disk_mem[ 9360] = 0;
disk_mem[ 9361] = 0;
disk_mem[ 9362] = 0;
disk_mem[ 9363] = 0;
disk_mem[ 9364] = 0;
disk_mem[ 9365] = 0;
disk_mem[ 9366] = 0;
disk_mem[ 9367] = 0;
disk_mem[ 9368] = 0;
disk_mem[ 9369] = 0;
disk_mem[ 9370] = 0;
disk_mem[ 9371] = 0;
disk_mem[ 9372] = 0;
disk_mem[ 9373] = 0;
disk_mem[ 9374] = 0;
disk_mem[ 9375] = 0;
disk_mem[ 9376] = 0;
disk_mem[ 9377] = 0;
disk_mem[ 9378] = 0;
disk_mem[ 9379] = 0;
disk_mem[ 9380] = 0;
disk_mem[ 9381] = 0;
disk_mem[ 9382] = 0;
disk_mem[ 9383] = 0;
disk_mem[ 9384] = 0;
disk_mem[ 9385] = 0;
disk_mem[ 9386] = 0;
disk_mem[ 9387] = 0;
disk_mem[ 9388] = 0;
disk_mem[ 9389] = 0;
disk_mem[ 9390] = 0;
disk_mem[ 9391] = 0;
disk_mem[ 9392] = 0;
disk_mem[ 9393] = 0;
disk_mem[ 9394] = 0;
disk_mem[ 9395] = 0;
disk_mem[ 9396] = 0;
disk_mem[ 9397] = 0;
disk_mem[ 9398] = 0;
disk_mem[ 9399] = 0;
disk_mem[ 9400] = 0;
disk_mem[ 9401] = 0;
disk_mem[ 9402] = 0;
disk_mem[ 9403] = 0;
disk_mem[ 9404] = 0;
disk_mem[ 9405] = 0;
disk_mem[ 9406] = 0;
disk_mem[ 9407] = 0;
disk_mem[ 9408] = 0;
disk_mem[ 9409] = 0;
disk_mem[ 9410] = 0;
disk_mem[ 9411] = 0;
disk_mem[ 9412] = 0;
disk_mem[ 9413] = 0;
disk_mem[ 9414] = 0;
disk_mem[ 9415] = 0;
disk_mem[ 9416] = 0;
disk_mem[ 9417] = 0;
disk_mem[ 9418] = 0;
disk_mem[ 9419] = 0;
disk_mem[ 9420] = 0;
disk_mem[ 9421] = 0;
disk_mem[ 9422] = 0;
disk_mem[ 9423] = 0;
disk_mem[ 9424] = 0;
disk_mem[ 9425] = 0;
disk_mem[ 9426] = 0;
disk_mem[ 9427] = 0;
disk_mem[ 9428] = 0;
disk_mem[ 9429] = 0;
disk_mem[ 9430] = 0;
disk_mem[ 9431] = 0;
disk_mem[ 9432] = 0;
disk_mem[ 9433] = 0;
disk_mem[ 9434] = 0;
disk_mem[ 9435] = 0;
disk_mem[ 9436] = 0;
disk_mem[ 9437] = 0;
disk_mem[ 9438] = 0;
disk_mem[ 9439] = 0;
disk_mem[ 9440] = 0;
disk_mem[ 9441] = 0;
disk_mem[ 9442] = 0;
disk_mem[ 9443] = 0;
disk_mem[ 9444] = 0;
disk_mem[ 9445] = 0;
disk_mem[ 9446] = 0;
disk_mem[ 9447] = 0;
disk_mem[ 9448] = 0;
disk_mem[ 9449] = 0;
disk_mem[ 9450] = 0;
disk_mem[ 9451] = 0;
disk_mem[ 9452] = 0;
disk_mem[ 9453] = 0;
disk_mem[ 9454] = 0;
disk_mem[ 9455] = 0;
disk_mem[ 9456] = 0;
disk_mem[ 9457] = 0;
disk_mem[ 9458] = 0;
disk_mem[ 9459] = 0;
disk_mem[ 9460] = 0;
disk_mem[ 9461] = 0;
disk_mem[ 9462] = 0;
disk_mem[ 9463] = 0;
disk_mem[ 9464] = 0;
disk_mem[ 9465] = 0;
disk_mem[ 9466] = 0;
disk_mem[ 9467] = 0;
disk_mem[ 9468] = 0;
disk_mem[ 9469] = 0;
disk_mem[ 9470] = 0;
disk_mem[ 9471] = 0;
disk_mem[ 9472] = 0;
disk_mem[ 9473] = 0;
disk_mem[ 9474] = 0;
disk_mem[ 9475] = 0;
disk_mem[ 9476] = 0;
disk_mem[ 9477] = 0;
disk_mem[ 9478] = 0;
disk_mem[ 9479] = 0;
disk_mem[ 9480] = 0;
disk_mem[ 9481] = 0;
disk_mem[ 9482] = 0;
disk_mem[ 9483] = 0;
disk_mem[ 9484] = 0;
disk_mem[ 9485] = 0;
disk_mem[ 9486] = 0;
disk_mem[ 9487] = 0;
disk_mem[ 9488] = 0;
disk_mem[ 9489] = 0;
disk_mem[ 9490] = 0;
disk_mem[ 9491] = 0;
disk_mem[ 9492] = 0;
disk_mem[ 9493] = 0;
disk_mem[ 9494] = 0;
disk_mem[ 9495] = 0;
disk_mem[ 9496] = 0;
disk_mem[ 9497] = 0;
disk_mem[ 9498] = 0;
disk_mem[ 9499] = 0;
disk_mem[ 9500] = 0;
disk_mem[ 9501] = 0;
disk_mem[ 9502] = 0;
disk_mem[ 9503] = 0;
disk_mem[ 9504] = 0;
disk_mem[ 9505] = 0;
disk_mem[ 9506] = 0;
disk_mem[ 9507] = 0;
disk_mem[ 9508] = 0;
disk_mem[ 9509] = 0;
disk_mem[ 9510] = 0;
disk_mem[ 9511] = 0;
disk_mem[ 9512] = 0;
disk_mem[ 9513] = 0;
disk_mem[ 9514] = 0;
disk_mem[ 9515] = 0;
disk_mem[ 9516] = 0;
disk_mem[ 9517] = 0;
disk_mem[ 9518] = 0;
disk_mem[ 9519] = 0;
disk_mem[ 9520] = 0;
disk_mem[ 9521] = 0;
disk_mem[ 9522] = 0;
disk_mem[ 9523] = 0;
disk_mem[ 9524] = 0;
disk_mem[ 9525] = 0;
disk_mem[ 9526] = 0;
disk_mem[ 9527] = 0;
disk_mem[ 9528] = 0;
disk_mem[ 9529] = 0;
disk_mem[ 9530] = 0;
disk_mem[ 9531] = 0;
disk_mem[ 9532] = 0;
disk_mem[ 9533] = 0;
disk_mem[ 9534] = 0;
disk_mem[ 9535] = 0;
disk_mem[ 9536] = 0;
disk_mem[ 9537] = 0;
disk_mem[ 9538] = 0;
disk_mem[ 9539] = 0;
disk_mem[ 9540] = 0;
disk_mem[ 9541] = 0;
disk_mem[ 9542] = 0;
disk_mem[ 9543] = 0;
disk_mem[ 9544] = 0;
disk_mem[ 9545] = 0;
disk_mem[ 9546] = 0;
disk_mem[ 9547] = 0;
disk_mem[ 9548] = 0;
disk_mem[ 9549] = 0;
disk_mem[ 9550] = 0;
disk_mem[ 9551] = 0;
disk_mem[ 9552] = 0;
disk_mem[ 9553] = 0;
disk_mem[ 9554] = 0;
disk_mem[ 9555] = 0;
disk_mem[ 9556] = 0;
disk_mem[ 9557] = 0;
disk_mem[ 9558] = 0;
disk_mem[ 9559] = 0;
disk_mem[ 9560] = 0;
disk_mem[ 9561] = 0;
disk_mem[ 9562] = 0;
disk_mem[ 9563] = 0;
disk_mem[ 9564] = 0;
disk_mem[ 9565] = 0;
disk_mem[ 9566] = 0;
disk_mem[ 9567] = 0;
disk_mem[ 9568] = 0;
disk_mem[ 9569] = 0;
disk_mem[ 9570] = 0;
disk_mem[ 9571] = 0;
disk_mem[ 9572] = 0;
disk_mem[ 9573] = 0;
disk_mem[ 9574] = 0;
disk_mem[ 9575] = 0;
disk_mem[ 9576] = 0;
disk_mem[ 9577] = 0;
disk_mem[ 9578] = 0;
disk_mem[ 9579] = 0;
disk_mem[ 9580] = 0;
disk_mem[ 9581] = 0;
disk_mem[ 9582] = 0;
disk_mem[ 9583] = 0;
disk_mem[ 9584] = 0;
disk_mem[ 9585] = 0;
disk_mem[ 9586] = 0;
disk_mem[ 9587] = 0;
disk_mem[ 9588] = 0;
disk_mem[ 9589] = 0;
disk_mem[ 9590] = 0;
disk_mem[ 9591] = 0;
disk_mem[ 9592] = 0;
disk_mem[ 9593] = 0;
disk_mem[ 9594] = 0;
disk_mem[ 9595] = 0;
disk_mem[ 9596] = 0;
disk_mem[ 9597] = 0;
disk_mem[ 9598] = 0;
disk_mem[ 9599] = 0;
disk_mem[ 9600] = 0;
disk_mem[ 9601] = 0;
disk_mem[ 9602] = 0;
disk_mem[ 9603] = 0;
disk_mem[ 9604] = 0;
disk_mem[ 9605] = 0;
disk_mem[ 9606] = 0;
disk_mem[ 9607] = 0;
disk_mem[ 9608] = 0;
disk_mem[ 9609] = 0;
disk_mem[ 9610] = 0;
disk_mem[ 9611] = 0;
disk_mem[ 9612] = 0;
disk_mem[ 9613] = 0;
disk_mem[ 9614] = 0;
disk_mem[ 9615] = 0;
disk_mem[ 9616] = 0;
disk_mem[ 9617] = 0;
disk_mem[ 9618] = 0;
disk_mem[ 9619] = 0;
disk_mem[ 9620] = 0;
disk_mem[ 9621] = 0;
disk_mem[ 9622] = 0;
disk_mem[ 9623] = 0;
disk_mem[ 9624] = 0;
disk_mem[ 9625] = 0;
disk_mem[ 9626] = 0;
disk_mem[ 9627] = 0;
disk_mem[ 9628] = 0;
disk_mem[ 9629] = 0;
disk_mem[ 9630] = 0;
disk_mem[ 9631] = 0;
disk_mem[ 9632] = 0;
disk_mem[ 9633] = 0;
disk_mem[ 9634] = 0;
disk_mem[ 9635] = 0;
disk_mem[ 9636] = 0;
disk_mem[ 9637] = 0;
disk_mem[ 9638] = 0;
disk_mem[ 9639] = 0;
disk_mem[ 9640] = 0;
disk_mem[ 9641] = 0;
disk_mem[ 9642] = 0;
disk_mem[ 9643] = 0;
disk_mem[ 9644] = 0;
disk_mem[ 9645] = 0;
disk_mem[ 9646] = 0;
disk_mem[ 9647] = 0;
disk_mem[ 9648] = 0;
disk_mem[ 9649] = 0;
disk_mem[ 9650] = 0;
disk_mem[ 9651] = 0;
disk_mem[ 9652] = 0;
disk_mem[ 9653] = 0;
disk_mem[ 9654] = 0;
disk_mem[ 9655] = 0;
disk_mem[ 9656] = 0;
disk_mem[ 9657] = 0;
disk_mem[ 9658] = 0;
disk_mem[ 9659] = 0;
disk_mem[ 9660] = 0;
disk_mem[ 9661] = 0;
disk_mem[ 9662] = 0;
disk_mem[ 9663] = 0;
disk_mem[ 9664] = 0;
disk_mem[ 9665] = 0;
disk_mem[ 9666] = 0;
disk_mem[ 9667] = 0;
disk_mem[ 9668] = 0;
disk_mem[ 9669] = 0;
disk_mem[ 9670] = 0;
disk_mem[ 9671] = 0;
disk_mem[ 9672] = 0;
disk_mem[ 9673] = 0;
disk_mem[ 9674] = 0;
disk_mem[ 9675] = 0;
disk_mem[ 9676] = 0;
disk_mem[ 9677] = 0;
disk_mem[ 9678] = 0;
disk_mem[ 9679] = 0;
disk_mem[ 9680] = 0;
disk_mem[ 9681] = 0;
disk_mem[ 9682] = 0;
disk_mem[ 9683] = 0;
disk_mem[ 9684] = 0;
disk_mem[ 9685] = 0;
disk_mem[ 9686] = 0;
disk_mem[ 9687] = 0;
disk_mem[ 9688] = 0;
disk_mem[ 9689] = 0;
disk_mem[ 9690] = 0;
disk_mem[ 9691] = 0;
disk_mem[ 9692] = 0;
disk_mem[ 9693] = 0;
disk_mem[ 9694] = 0;
disk_mem[ 9695] = 0;
disk_mem[ 9696] = 0;
disk_mem[ 9697] = 0;
disk_mem[ 9698] = 0;
disk_mem[ 9699] = 0;
disk_mem[ 9700] = 0;
disk_mem[ 9701] = 0;
disk_mem[ 9702] = 0;
disk_mem[ 9703] = 0;
disk_mem[ 9704] = 0;
disk_mem[ 9705] = 0;
disk_mem[ 9706] = 0;
disk_mem[ 9707] = 0;
disk_mem[ 9708] = 0;
disk_mem[ 9709] = 0;
disk_mem[ 9710] = 0;
disk_mem[ 9711] = 0;
disk_mem[ 9712] = 0;
disk_mem[ 9713] = 0;
disk_mem[ 9714] = 0;
disk_mem[ 9715] = 0;
disk_mem[ 9716] = 0;
disk_mem[ 9717] = 0;
disk_mem[ 9718] = 0;
disk_mem[ 9719] = 0;
disk_mem[ 9720] = 0;
disk_mem[ 9721] = 0;
disk_mem[ 9722] = 0;
disk_mem[ 9723] = 0;
disk_mem[ 9724] = 0;
disk_mem[ 9725] = 0;
disk_mem[ 9726] = 0;
disk_mem[ 9727] = 0;
disk_mem[ 9728] = 0;
disk_mem[ 9729] = 0;
disk_mem[ 9730] = 0;
disk_mem[ 9731] = 0;
disk_mem[ 9732] = 0;
disk_mem[ 9733] = 0;
disk_mem[ 9734] = 0;
disk_mem[ 9735] = 0;
disk_mem[ 9736] = 0;
disk_mem[ 9737] = 0;
disk_mem[ 9738] = 0;
disk_mem[ 9739] = 0;
disk_mem[ 9740] = 0;
disk_mem[ 9741] = 0;
disk_mem[ 9742] = 0;
disk_mem[ 9743] = 0;
disk_mem[ 9744] = 0;
disk_mem[ 9745] = 0;
disk_mem[ 9746] = 0;
disk_mem[ 9747] = 0;
disk_mem[ 9748] = 0;
disk_mem[ 9749] = 0;
disk_mem[ 9750] = 0;
disk_mem[ 9751] = 0;
disk_mem[ 9752] = 0;
disk_mem[ 9753] = 0;
disk_mem[ 9754] = 0;
disk_mem[ 9755] = 0;
disk_mem[ 9756] = 0;
disk_mem[ 9757] = 0;
disk_mem[ 9758] = 0;
disk_mem[ 9759] = 0;
disk_mem[ 9760] = 0;
disk_mem[ 9761] = 0;
disk_mem[ 9762] = 0;
disk_mem[ 9763] = 0;
disk_mem[ 9764] = 0;
disk_mem[ 9765] = 0;
disk_mem[ 9766] = 0;
disk_mem[ 9767] = 0;
disk_mem[ 9768] = 0;
disk_mem[ 9769] = 0;
disk_mem[ 9770] = 0;
disk_mem[ 9771] = 0;
disk_mem[ 9772] = 0;
disk_mem[ 9773] = 0;
disk_mem[ 9774] = 0;
disk_mem[ 9775] = 0;
disk_mem[ 9776] = 0;
disk_mem[ 9777] = 0;
disk_mem[ 9778] = 0;
disk_mem[ 9779] = 0;
disk_mem[ 9780] = 0;
disk_mem[ 9781] = 0;
disk_mem[ 9782] = 0;
disk_mem[ 9783] = 0;
disk_mem[ 9784] = 0;
disk_mem[ 9785] = 0;
disk_mem[ 9786] = 0;
disk_mem[ 9787] = 0;
disk_mem[ 9788] = 0;
disk_mem[ 9789] = 0;
disk_mem[ 9790] = 0;
disk_mem[ 9791] = 0;
disk_mem[ 9792] = 0;
disk_mem[ 9793] = 0;
disk_mem[ 9794] = 0;
disk_mem[ 9795] = 0;
disk_mem[ 9796] = 0;
disk_mem[ 9797] = 0;
disk_mem[ 9798] = 0;
disk_mem[ 9799] = 0;
disk_mem[ 9800] = 0;
disk_mem[ 9801] = 0;
disk_mem[ 9802] = 0;
disk_mem[ 9803] = 0;
disk_mem[ 9804] = 0;
disk_mem[ 9805] = 0;
disk_mem[ 9806] = 0;
disk_mem[ 9807] = 0;
disk_mem[ 9808] = 0;
disk_mem[ 9809] = 0;
disk_mem[ 9810] = 0;
disk_mem[ 9811] = 0;
disk_mem[ 9812] = 0;
disk_mem[ 9813] = 0;
disk_mem[ 9814] = 0;
disk_mem[ 9815] = 0;
disk_mem[ 9816] = 0;
disk_mem[ 9817] = 0;
disk_mem[ 9818] = 0;
disk_mem[ 9819] = 0;
disk_mem[ 9820] = 0;
disk_mem[ 9821] = 0;
disk_mem[ 9822] = 0;
disk_mem[ 9823] = 0;
disk_mem[ 9824] = 0;
disk_mem[ 9825] = 0;
disk_mem[ 9826] = 0;
disk_mem[ 9827] = 0;
disk_mem[ 9828] = 0;
disk_mem[ 9829] = 0;
disk_mem[ 9830] = 0;
disk_mem[ 9831] = 0;
disk_mem[ 9832] = 0;
disk_mem[ 9833] = 0;
disk_mem[ 9834] = 0;
disk_mem[ 9835] = 0;
disk_mem[ 9836] = 0;
disk_mem[ 9837] = 0;
disk_mem[ 9838] = 0;
disk_mem[ 9839] = 0;
disk_mem[ 9840] = 0;
disk_mem[ 9841] = 0;
disk_mem[ 9842] = 0;
disk_mem[ 9843] = 0;
disk_mem[ 9844] = 0;
disk_mem[ 9845] = 0;
disk_mem[ 9846] = 0;
disk_mem[ 9847] = 0;
disk_mem[ 9848] = 0;
disk_mem[ 9849] = 0;
disk_mem[ 9850] = 0;
disk_mem[ 9851] = 0;
disk_mem[ 9852] = 0;
disk_mem[ 9853] = 0;
disk_mem[ 9854] = 0;
disk_mem[ 9855] = 0;
disk_mem[ 9856] = 0;
disk_mem[ 9857] = 0;
disk_mem[ 9858] = 0;
disk_mem[ 9859] = 0;
disk_mem[ 9860] = 0;
disk_mem[ 9861] = 0;
disk_mem[ 9862] = 0;
disk_mem[ 9863] = 0;
disk_mem[ 9864] = 0;
disk_mem[ 9865] = 0;
disk_mem[ 9866] = 0;
disk_mem[ 9867] = 0;
disk_mem[ 9868] = 0;
disk_mem[ 9869] = 0;
disk_mem[ 9870] = 0;
disk_mem[ 9871] = 0;
disk_mem[ 9872] = 0;
disk_mem[ 9873] = 0;
disk_mem[ 9874] = 0;
disk_mem[ 9875] = 0;
disk_mem[ 9876] = 0;
disk_mem[ 9877] = 0;
disk_mem[ 9878] = 0;
disk_mem[ 9879] = 0;
disk_mem[ 9880] = 0;
disk_mem[ 9881] = 0;
disk_mem[ 9882] = 0;
disk_mem[ 9883] = 0;
disk_mem[ 9884] = 0;
disk_mem[ 9885] = 0;
disk_mem[ 9886] = 0;
disk_mem[ 9887] = 0;
disk_mem[ 9888] = 0;
disk_mem[ 9889] = 0;
disk_mem[ 9890] = 0;
disk_mem[ 9891] = 0;
disk_mem[ 9892] = 0;
disk_mem[ 9893] = 0;
disk_mem[ 9894] = 0;
disk_mem[ 9895] = 0;
disk_mem[ 9896] = 0;
disk_mem[ 9897] = 0;
disk_mem[ 9898] = 0;
disk_mem[ 9899] = 0;
disk_mem[ 9900] = 0;
disk_mem[ 9901] = 0;
disk_mem[ 9902] = 0;
disk_mem[ 9903] = 0;
disk_mem[ 9904] = 0;
disk_mem[ 9905] = 0;
disk_mem[ 9906] = 0;
disk_mem[ 9907] = 0;
disk_mem[ 9908] = 0;
disk_mem[ 9909] = 0;
disk_mem[ 9910] = 0;
disk_mem[ 9911] = 0;
disk_mem[ 9912] = 0;
disk_mem[ 9913] = 0;
disk_mem[ 9914] = 0;
disk_mem[ 9915] = 0;
disk_mem[ 9916] = 0;
disk_mem[ 9917] = 0;
disk_mem[ 9918] = 0;
disk_mem[ 9919] = 0;
disk_mem[ 9920] = 0;
disk_mem[ 9921] = 0;
disk_mem[ 9922] = 0;
disk_mem[ 9923] = 0;
disk_mem[ 9924] = 0;
disk_mem[ 9925] = 0;
disk_mem[ 9926] = 0;
disk_mem[ 9927] = 0;
disk_mem[ 9928] = 0;
disk_mem[ 9929] = 0;
disk_mem[ 9930] = 0;
disk_mem[ 9931] = 0;
disk_mem[ 9932] = 0;
disk_mem[ 9933] = 0;
disk_mem[ 9934] = 0;
disk_mem[ 9935] = 0;
disk_mem[ 9936] = 0;
disk_mem[ 9937] = 0;
disk_mem[ 9938] = 0;
disk_mem[ 9939] = 0;
disk_mem[ 9940] = 0;
disk_mem[ 9941] = 0;
disk_mem[ 9942] = 0;
disk_mem[ 9943] = 0;
disk_mem[ 9944] = 0;
disk_mem[ 9945] = 0;
disk_mem[ 9946] = 0;
disk_mem[ 9947] = 0;
disk_mem[ 9948] = 0;
disk_mem[ 9949] = 0;
disk_mem[ 9950] = 0;
disk_mem[ 9951] = 0;
disk_mem[ 9952] = 0;
disk_mem[ 9953] = 0;
disk_mem[ 9954] = 0;
disk_mem[ 9955] = 0;
disk_mem[ 9956] = 0;
disk_mem[ 9957] = 0;
disk_mem[ 9958] = 0;
disk_mem[ 9959] = 0;
disk_mem[ 9960] = 0;
disk_mem[ 9961] = 0;
disk_mem[ 9962] = 0;
disk_mem[ 9963] = 0;
disk_mem[ 9964] = 0;
disk_mem[ 9965] = 0;
disk_mem[ 9966] = 0;
disk_mem[ 9967] = 0;
disk_mem[ 9968] = 0;
disk_mem[ 9969] = 0;
disk_mem[ 9970] = 0;
disk_mem[ 9971] = 0;
disk_mem[ 9972] = 0;
disk_mem[ 9973] = 0;
disk_mem[ 9974] = 0;
disk_mem[ 9975] = 0;
disk_mem[ 9976] = 0;
disk_mem[ 9977] = 0;
disk_mem[ 9978] = 0;
disk_mem[ 9979] = 0;
disk_mem[ 9980] = 0;
disk_mem[ 9981] = 0;
disk_mem[ 9982] = 0;
disk_mem[ 9983] = 0;
disk_mem[ 9984] = 0;
disk_mem[ 9985] = 0;
disk_mem[ 9986] = 0;
disk_mem[ 9987] = 0;
disk_mem[ 9988] = 0;
disk_mem[ 9989] = 0;
disk_mem[ 9990] = 0;
disk_mem[ 9991] = 0;
disk_mem[ 9992] = 0;
disk_mem[ 9993] = 0;
disk_mem[ 9994] = 0;
disk_mem[ 9995] = 0;
disk_mem[ 9996] = 0;
disk_mem[ 9997] = 0;
disk_mem[ 9998] = 0;
disk_mem[ 9999] = 0;
disk_mem[10000] = 0;
disk_mem[10001] = 0;
disk_mem[10002] = 0;
disk_mem[10003] = 0;
disk_mem[10004] = 0;
disk_mem[10005] = 0;
disk_mem[10006] = 0;
disk_mem[10007] = 0;
disk_mem[10008] = 0;
disk_mem[10009] = 0;
disk_mem[10010] = 0;
disk_mem[10011] = 0;
disk_mem[10012] = 0;
disk_mem[10013] = 0;
disk_mem[10014] = 0;
disk_mem[10015] = 0;
disk_mem[10016] = 0;
disk_mem[10017] = 0;
disk_mem[10018] = 0;
disk_mem[10019] = 0;
disk_mem[10020] = 0;
disk_mem[10021] = 0;
disk_mem[10022] = 0;
disk_mem[10023] = 0;
disk_mem[10024] = 0;
disk_mem[10025] = 0;
disk_mem[10026] = 0;
disk_mem[10027] = 0;
disk_mem[10028] = 0;
disk_mem[10029] = 0;
disk_mem[10030] = 0;
disk_mem[10031] = 0;
disk_mem[10032] = 0;
disk_mem[10033] = 0;
disk_mem[10034] = 0;
disk_mem[10035] = 0;
disk_mem[10036] = 0;
disk_mem[10037] = 0;
disk_mem[10038] = 0;
disk_mem[10039] = 0;
disk_mem[10040] = 0;
disk_mem[10041] = 0;
disk_mem[10042] = 0;
disk_mem[10043] = 0;
disk_mem[10044] = 0;
disk_mem[10045] = 0;
disk_mem[10046] = 0;
disk_mem[10047] = 0;
disk_mem[10048] = 0;
disk_mem[10049] = 0;
disk_mem[10050] = 0;
disk_mem[10051] = 0;
disk_mem[10052] = 0;
disk_mem[10053] = 0;
disk_mem[10054] = 0;
disk_mem[10055] = 0;
disk_mem[10056] = 0;
disk_mem[10057] = 0;
disk_mem[10058] = 0;
disk_mem[10059] = 0;
disk_mem[10060] = 0;
disk_mem[10061] = 0;
disk_mem[10062] = 0;
disk_mem[10063] = 0;
disk_mem[10064] = 0;
disk_mem[10065] = 0;
disk_mem[10066] = 0;
disk_mem[10067] = 0;
disk_mem[10068] = 0;
disk_mem[10069] = 0;
disk_mem[10070] = 0;
disk_mem[10071] = 0;
disk_mem[10072] = 0;
disk_mem[10073] = 0;
disk_mem[10074] = 0;
disk_mem[10075] = 0;
disk_mem[10076] = 0;
disk_mem[10077] = 0;
disk_mem[10078] = 0;
disk_mem[10079] = 0;
disk_mem[10080] = 0;
disk_mem[10081] = 0;
disk_mem[10082] = 0;
disk_mem[10083] = 0;
disk_mem[10084] = 0;
disk_mem[10085] = 0;
disk_mem[10086] = 0;
disk_mem[10087] = 0;
disk_mem[10088] = 0;
disk_mem[10089] = 0;
disk_mem[10090] = 0;
disk_mem[10091] = 0;
disk_mem[10092] = 0;
disk_mem[10093] = 0;
disk_mem[10094] = 0;
disk_mem[10095] = 0;
disk_mem[10096] = 0;
disk_mem[10097] = 0;
disk_mem[10098] = 0;
disk_mem[10099] = 0;
disk_mem[10100] = 0;
disk_mem[10101] = 0;
disk_mem[10102] = 0;
disk_mem[10103] = 0;
disk_mem[10104] = 0;
disk_mem[10105] = 0;
disk_mem[10106] = 0;
disk_mem[10107] = 0;
disk_mem[10108] = 0;
disk_mem[10109] = 0;
disk_mem[10110] = 0;
disk_mem[10111] = 0;
disk_mem[10112] = 0;
disk_mem[10113] = 0;
disk_mem[10114] = 0;
disk_mem[10115] = 0;
disk_mem[10116] = 0;
disk_mem[10117] = 0;
disk_mem[10118] = 0;
disk_mem[10119] = 0;
disk_mem[10120] = 0;
disk_mem[10121] = 0;
disk_mem[10122] = 0;
disk_mem[10123] = 0;
disk_mem[10124] = 0;
disk_mem[10125] = 0;
disk_mem[10126] = 0;
disk_mem[10127] = 0;
disk_mem[10128] = 0;
disk_mem[10129] = 0;
disk_mem[10130] = 0;
disk_mem[10131] = 0;
disk_mem[10132] = 0;
disk_mem[10133] = 0;
disk_mem[10134] = 0;
disk_mem[10135] = 0;
disk_mem[10136] = 0;
disk_mem[10137] = 0;
disk_mem[10138] = 0;
disk_mem[10139] = 0;
disk_mem[10140] = 0;
disk_mem[10141] = 0;
disk_mem[10142] = 0;
disk_mem[10143] = 0;
disk_mem[10144] = 0;
disk_mem[10145] = 0;
disk_mem[10146] = 0;
disk_mem[10147] = 0;
disk_mem[10148] = 0;
disk_mem[10149] = 0;
disk_mem[10150] = 0;
disk_mem[10151] = 0;
disk_mem[10152] = 0;
disk_mem[10153] = 0;
disk_mem[10154] = 0;
disk_mem[10155] = 0;
disk_mem[10156] = 0;
disk_mem[10157] = 0;
disk_mem[10158] = 0;
disk_mem[10159] = 0;
disk_mem[10160] = 0;
disk_mem[10161] = 0;
disk_mem[10162] = 0;
disk_mem[10163] = 0;
disk_mem[10164] = 0;
disk_mem[10165] = 0;
disk_mem[10166] = 0;
disk_mem[10167] = 0;
disk_mem[10168] = 0;
disk_mem[10169] = 0;
disk_mem[10170] = 0;
disk_mem[10171] = 0;
disk_mem[10172] = 0;
disk_mem[10173] = 0;
disk_mem[10174] = 0;
disk_mem[10175] = 0;
disk_mem[10176] = 0;
disk_mem[10177] = 0;
disk_mem[10178] = 0;
disk_mem[10179] = 0;
disk_mem[10180] = 0;
disk_mem[10181] = 0;
disk_mem[10182] = 0;
disk_mem[10183] = 0;
disk_mem[10184] = 0;
disk_mem[10185] = 0;
disk_mem[10186] = 0;
disk_mem[10187] = 0;
disk_mem[10188] = 0;
disk_mem[10189] = 0;
disk_mem[10190] = 0;
disk_mem[10191] = 0;
disk_mem[10192] = 0;
disk_mem[10193] = 0;
disk_mem[10194] = 0;
disk_mem[10195] = 0;
disk_mem[10196] = 0;
disk_mem[10197] = 0;
disk_mem[10198] = 0;
disk_mem[10199] = 0;
disk_mem[10200] = 0;
disk_mem[10201] = 0;
disk_mem[10202] = 0;
disk_mem[10203] = 0;
disk_mem[10204] = 0;
disk_mem[10205] = 0;
disk_mem[10206] = 0;
disk_mem[10207] = 0;
disk_mem[10208] = 0;
disk_mem[10209] = 0;
disk_mem[10210] = 0;
disk_mem[10211] = 0;
disk_mem[10212] = 0;
disk_mem[10213] = 0;
disk_mem[10214] = 0;
disk_mem[10215] = 0;
disk_mem[10216] = 0;
disk_mem[10217] = 0;
disk_mem[10218] = 0;
disk_mem[10219] = 0;
disk_mem[10220] = 0;
disk_mem[10221] = 0;
disk_mem[10222] = 0;
disk_mem[10223] = 0;
disk_mem[10224] = 0;
disk_mem[10225] = 0;
disk_mem[10226] = 0;
disk_mem[10227] = 0;
disk_mem[10228] = 0;
disk_mem[10229] = 0;
disk_mem[10230] = 0;
disk_mem[10231] = 0;
disk_mem[10232] = 0;
disk_mem[10233] = 0;
disk_mem[10234] = 0;
disk_mem[10235] = 0;
disk_mem[10236] = 0;
disk_mem[10237] = 0;
disk_mem[10238] = 0;
disk_mem[10239] = 0;
disk_mem[10240] = 0;
disk_mem[10241] = 0;
disk_mem[10242] = 0;
disk_mem[10243] = 0;
disk_mem[10244] = 0;
disk_mem[10245] = 0;
disk_mem[10246] = 0;
disk_mem[10247] = 0;
disk_mem[10248] = 0;
disk_mem[10249] = 0;
disk_mem[10250] = 0;
disk_mem[10251] = 0;
disk_mem[10252] = 0;
disk_mem[10253] = 0;
disk_mem[10254] = 0;
disk_mem[10255] = 0;
disk_mem[10256] = 0;
disk_mem[10257] = 0;
disk_mem[10258] = 0;
disk_mem[10259] = 0;
disk_mem[10260] = 0;
disk_mem[10261] = 0;
disk_mem[10262] = 0;
disk_mem[10263] = 0;
disk_mem[10264] = 0;
disk_mem[10265] = 0;
disk_mem[10266] = 0;
disk_mem[10267] = 0;
disk_mem[10268] = 0;
disk_mem[10269] = 0;
disk_mem[10270] = 0;
disk_mem[10271] = 0;
disk_mem[10272] = 0;
disk_mem[10273] = 0;
disk_mem[10274] = 0;
disk_mem[10275] = 0;
disk_mem[10276] = 0;
disk_mem[10277] = 0;
disk_mem[10278] = 0;
disk_mem[10279] = 0;
disk_mem[10280] = 0;
disk_mem[10281] = 0;
disk_mem[10282] = 0;
disk_mem[10283] = 0;
disk_mem[10284] = 0;
disk_mem[10285] = 0;
disk_mem[10286] = 0;
disk_mem[10287] = 0;
disk_mem[10288] = 0;
disk_mem[10289] = 0;
disk_mem[10290] = 0;
disk_mem[10291] = 0;
disk_mem[10292] = 0;
disk_mem[10293] = 0;
disk_mem[10294] = 0;
disk_mem[10295] = 0;
disk_mem[10296] = 0;
disk_mem[10297] = 0;
disk_mem[10298] = 0;
disk_mem[10299] = 0;
disk_mem[10300] = 0;
disk_mem[10301] = 0;
disk_mem[10302] = 0;
disk_mem[10303] = 0;
disk_mem[10304] = 0;
disk_mem[10305] = 0;
disk_mem[10306] = 0;
disk_mem[10307] = 0;
disk_mem[10308] = 0;
disk_mem[10309] = 0;
disk_mem[10310] = 0;
disk_mem[10311] = 0;
disk_mem[10312] = 0;
disk_mem[10313] = 0;
disk_mem[10314] = 0;
disk_mem[10315] = 0;
disk_mem[10316] = 0;
disk_mem[10317] = 0;
disk_mem[10318] = 0;
disk_mem[10319] = 0;
disk_mem[10320] = 0;
disk_mem[10321] = 0;
disk_mem[10322] = 0;
disk_mem[10323] = 0;
disk_mem[10324] = 0;
disk_mem[10325] = 0;
disk_mem[10326] = 0;
disk_mem[10327] = 0;
disk_mem[10328] = 0;
disk_mem[10329] = 0;
disk_mem[10330] = 0;
disk_mem[10331] = 0;
disk_mem[10332] = 0;
disk_mem[10333] = 0;
disk_mem[10334] = 0;
disk_mem[10335] = 0;
disk_mem[10336] = 0;
disk_mem[10337] = 0;
disk_mem[10338] = 0;
disk_mem[10339] = 0;
disk_mem[10340] = 0;
disk_mem[10341] = 0;
disk_mem[10342] = 0;
disk_mem[10343] = 0;
disk_mem[10344] = 0;
disk_mem[10345] = 0;
disk_mem[10346] = 0;
disk_mem[10347] = 0;
disk_mem[10348] = 0;
disk_mem[10349] = 0;
disk_mem[10350] = 0;
disk_mem[10351] = 0;
disk_mem[10352] = 0;
disk_mem[10353] = 0;
disk_mem[10354] = 0;
disk_mem[10355] = 0;
disk_mem[10356] = 0;
disk_mem[10357] = 0;
disk_mem[10358] = 0;
disk_mem[10359] = 0;
disk_mem[10360] = 0;
disk_mem[10361] = 0;
disk_mem[10362] = 0;
disk_mem[10363] = 0;
disk_mem[10364] = 0;
disk_mem[10365] = 0;
disk_mem[10366] = 0;
disk_mem[10367] = 0;
disk_mem[10368] = 0;
disk_mem[10369] = 0;
disk_mem[10370] = 0;
disk_mem[10371] = 0;
disk_mem[10372] = 0;
disk_mem[10373] = 0;
disk_mem[10374] = 0;
disk_mem[10375] = 0;
disk_mem[10376] = 0;
disk_mem[10377] = 0;
disk_mem[10378] = 0;
disk_mem[10379] = 0;
disk_mem[10380] = 0;
disk_mem[10381] = 0;
disk_mem[10382] = 0;
disk_mem[10383] = 0;
disk_mem[10384] = 0;
disk_mem[10385] = 0;
disk_mem[10386] = 0;
disk_mem[10387] = 0;
disk_mem[10388] = 0;
disk_mem[10389] = 0;
disk_mem[10390] = 0;
disk_mem[10391] = 0;
disk_mem[10392] = 0;
disk_mem[10393] = 0;
disk_mem[10394] = 0;
disk_mem[10395] = 0;
disk_mem[10396] = 0;
disk_mem[10397] = 0;
disk_mem[10398] = 0;
disk_mem[10399] = 0;
disk_mem[10400] = 0;
disk_mem[10401] = 0;
disk_mem[10402] = 0;
disk_mem[10403] = 0;
disk_mem[10404] = 0;
disk_mem[10405] = 0;
disk_mem[10406] = 0;
disk_mem[10407] = 0;
disk_mem[10408] = 0;
disk_mem[10409] = 0;
disk_mem[10410] = 0;
disk_mem[10411] = 0;
disk_mem[10412] = 0;
disk_mem[10413] = 0;
disk_mem[10414] = 0;
disk_mem[10415] = 0;
disk_mem[10416] = 0;
disk_mem[10417] = 0;
disk_mem[10418] = 0;
disk_mem[10419] = 0;
disk_mem[10420] = 0;
disk_mem[10421] = 0;
disk_mem[10422] = 0;
disk_mem[10423] = 0;
disk_mem[10424] = 0;
disk_mem[10425] = 0;
disk_mem[10426] = 0;
disk_mem[10427] = 0;
disk_mem[10428] = 0;
disk_mem[10429] = 0;
disk_mem[10430] = 0;
disk_mem[10431] = 0;
disk_mem[10432] = 0;
disk_mem[10433] = 0;
disk_mem[10434] = 0;
disk_mem[10435] = 0;
disk_mem[10436] = 0;
disk_mem[10437] = 0;
disk_mem[10438] = 0;
disk_mem[10439] = 0;
disk_mem[10440] = 0;
disk_mem[10441] = 0;
disk_mem[10442] = 0;
disk_mem[10443] = 0;
disk_mem[10444] = 0;
disk_mem[10445] = 0;
disk_mem[10446] = 0;
disk_mem[10447] = 0;
disk_mem[10448] = 0;
disk_mem[10449] = 0;
disk_mem[10450] = 0;
disk_mem[10451] = 0;
disk_mem[10452] = 0;
disk_mem[10453] = 0;
disk_mem[10454] = 0;
disk_mem[10455] = 0;
disk_mem[10456] = 0;
disk_mem[10457] = 0;
disk_mem[10458] = 0;
disk_mem[10459] = 0;
disk_mem[10460] = 0;
disk_mem[10461] = 0;
disk_mem[10462] = 0;
disk_mem[10463] = 0;
disk_mem[10464] = 0;
disk_mem[10465] = 0;
disk_mem[10466] = 0;
disk_mem[10467] = 0;
disk_mem[10468] = 0;
disk_mem[10469] = 0;
disk_mem[10470] = 0;
disk_mem[10471] = 0;
disk_mem[10472] = 0;
disk_mem[10473] = 0;
disk_mem[10474] = 0;
disk_mem[10475] = 0;
disk_mem[10476] = 0;
disk_mem[10477] = 0;
disk_mem[10478] = 0;
disk_mem[10479] = 0;
disk_mem[10480] = 0;
disk_mem[10481] = 0;
disk_mem[10482] = 0;
disk_mem[10483] = 0;
disk_mem[10484] = 0;
disk_mem[10485] = 0;
disk_mem[10486] = 0;
disk_mem[10487] = 0;
disk_mem[10488] = 0;
disk_mem[10489] = 0;
disk_mem[10490] = 0;
disk_mem[10491] = 0;
disk_mem[10492] = 0;
disk_mem[10493] = 0;
disk_mem[10494] = 0;
disk_mem[10495] = 0;
disk_mem[10496] = 0;
disk_mem[10497] = 0;
disk_mem[10498] = 0;
disk_mem[10499] = 0;
disk_mem[10500] = 0;
disk_mem[10501] = 0;
disk_mem[10502] = 0;
disk_mem[10503] = 0;
disk_mem[10504] = 0;
disk_mem[10505] = 0;
disk_mem[10506] = 0;
disk_mem[10507] = 0;
disk_mem[10508] = 0;
disk_mem[10509] = 0;
disk_mem[10510] = 0;
disk_mem[10511] = 0;
disk_mem[10512] = 0;
disk_mem[10513] = 0;
disk_mem[10514] = 0;
disk_mem[10515] = 0;
disk_mem[10516] = 0;
disk_mem[10517] = 0;
disk_mem[10518] = 0;
disk_mem[10519] = 0;
disk_mem[10520] = 0;
disk_mem[10521] = 0;
disk_mem[10522] = 0;
disk_mem[10523] = 0;
disk_mem[10524] = 0;
disk_mem[10525] = 0;
disk_mem[10526] = 0;
disk_mem[10527] = 0;
disk_mem[10528] = 0;
disk_mem[10529] = 0;
disk_mem[10530] = 0;
disk_mem[10531] = 0;
disk_mem[10532] = 0;
disk_mem[10533] = 0;
disk_mem[10534] = 0;
disk_mem[10535] = 0;
disk_mem[10536] = 0;
disk_mem[10537] = 0;
disk_mem[10538] = 0;
disk_mem[10539] = 0;
disk_mem[10540] = 0;
disk_mem[10541] = 0;
disk_mem[10542] = 0;
disk_mem[10543] = 0;
disk_mem[10544] = 0;
disk_mem[10545] = 0;
disk_mem[10546] = 0;
disk_mem[10547] = 0;
disk_mem[10548] = 0;
disk_mem[10549] = 0;
disk_mem[10550] = 0;
disk_mem[10551] = 0;
disk_mem[10552] = 0;
disk_mem[10553] = 0;
disk_mem[10554] = 0;
disk_mem[10555] = 0;
disk_mem[10556] = 0;
disk_mem[10557] = 0;
disk_mem[10558] = 0;
disk_mem[10559] = 0;
disk_mem[10560] = 0;
disk_mem[10561] = 0;
disk_mem[10562] = 0;
disk_mem[10563] = 0;
disk_mem[10564] = 0;
disk_mem[10565] = 0;
disk_mem[10566] = 0;
disk_mem[10567] = 0;
disk_mem[10568] = 0;
disk_mem[10569] = 0;
disk_mem[10570] = 0;
disk_mem[10571] = 0;
disk_mem[10572] = 0;
disk_mem[10573] = 0;
disk_mem[10574] = 0;
disk_mem[10575] = 0;
disk_mem[10576] = 0;
disk_mem[10577] = 0;
disk_mem[10578] = 0;
disk_mem[10579] = 0;
disk_mem[10580] = 0;
disk_mem[10581] = 0;
disk_mem[10582] = 0;
disk_mem[10583] = 0;
disk_mem[10584] = 0;
disk_mem[10585] = 0;
disk_mem[10586] = 0;
disk_mem[10587] = 0;
disk_mem[10588] = 0;
disk_mem[10589] = 0;
disk_mem[10590] = 0;
disk_mem[10591] = 0;
disk_mem[10592] = 0;
disk_mem[10593] = 0;
disk_mem[10594] = 0;
disk_mem[10595] = 0;
disk_mem[10596] = 0;
disk_mem[10597] = 0;
disk_mem[10598] = 0;
disk_mem[10599] = 0;
disk_mem[10600] = 0;
disk_mem[10601] = 0;
disk_mem[10602] = 0;
disk_mem[10603] = 0;
disk_mem[10604] = 0;
disk_mem[10605] = 0;
disk_mem[10606] = 0;
disk_mem[10607] = 0;
disk_mem[10608] = 0;
disk_mem[10609] = 0;
disk_mem[10610] = 0;
disk_mem[10611] = 0;
disk_mem[10612] = 0;
disk_mem[10613] = 0;
disk_mem[10614] = 0;
disk_mem[10615] = 0;
disk_mem[10616] = 0;
disk_mem[10617] = 0;
disk_mem[10618] = 0;
disk_mem[10619] = 0;
disk_mem[10620] = 0;
disk_mem[10621] = 0;
disk_mem[10622] = 0;
disk_mem[10623] = 0;
disk_mem[10624] = 0;
disk_mem[10625] = 0;
disk_mem[10626] = 0;
disk_mem[10627] = 0;
disk_mem[10628] = 0;
disk_mem[10629] = 0;
disk_mem[10630] = 0;
disk_mem[10631] = 0;
disk_mem[10632] = 0;
disk_mem[10633] = 0;
disk_mem[10634] = 0;
disk_mem[10635] = 0;
disk_mem[10636] = 0;
disk_mem[10637] = 0;
disk_mem[10638] = 0;
disk_mem[10639] = 0;
disk_mem[10640] = 0;
disk_mem[10641] = 0;
disk_mem[10642] = 0;
disk_mem[10643] = 0;
disk_mem[10644] = 0;
disk_mem[10645] = 0;
disk_mem[10646] = 0;
disk_mem[10647] = 0;
disk_mem[10648] = 0;
disk_mem[10649] = 0;
disk_mem[10650] = 0;
disk_mem[10651] = 0;
disk_mem[10652] = 0;
disk_mem[10653] = 0;
disk_mem[10654] = 0;
disk_mem[10655] = 0;
disk_mem[10656] = 0;
disk_mem[10657] = 0;
disk_mem[10658] = 0;
disk_mem[10659] = 0;
disk_mem[10660] = 0;
disk_mem[10661] = 0;
disk_mem[10662] = 0;
disk_mem[10663] = 0;
disk_mem[10664] = 0;
disk_mem[10665] = 0;
disk_mem[10666] = 0;
disk_mem[10667] = 0;
disk_mem[10668] = 0;
disk_mem[10669] = 0;
disk_mem[10670] = 0;
disk_mem[10671] = 0;
disk_mem[10672] = 0;
disk_mem[10673] = 0;
disk_mem[10674] = 0;
disk_mem[10675] = 0;
disk_mem[10676] = 0;
disk_mem[10677] = 0;
disk_mem[10678] = 0;
disk_mem[10679] = 0;
disk_mem[10680] = 0;
disk_mem[10681] = 0;
disk_mem[10682] = 0;
disk_mem[10683] = 0;
disk_mem[10684] = 0;
disk_mem[10685] = 0;
disk_mem[10686] = 0;
disk_mem[10687] = 0;
disk_mem[10688] = 0;
disk_mem[10689] = 0;
disk_mem[10690] = 0;
disk_mem[10691] = 0;
disk_mem[10692] = 0;
disk_mem[10693] = 0;
disk_mem[10694] = 0;
disk_mem[10695] = 0;
disk_mem[10696] = 0;
disk_mem[10697] = 0;
disk_mem[10698] = 0;
disk_mem[10699] = 0;
disk_mem[10700] = 0;
disk_mem[10701] = 0;
disk_mem[10702] = 0;
disk_mem[10703] = 0;
disk_mem[10704] = 0;
disk_mem[10705] = 0;
disk_mem[10706] = 0;
disk_mem[10707] = 0;
disk_mem[10708] = 0;
disk_mem[10709] = 0;
disk_mem[10710] = 0;
disk_mem[10711] = 0;
disk_mem[10712] = 0;
disk_mem[10713] = 0;
disk_mem[10714] = 0;
disk_mem[10715] = 0;
disk_mem[10716] = 0;
disk_mem[10717] = 0;
disk_mem[10718] = 0;
disk_mem[10719] = 0;
disk_mem[10720] = 0;
disk_mem[10721] = 0;
disk_mem[10722] = 0;
disk_mem[10723] = 0;
disk_mem[10724] = 0;
disk_mem[10725] = 0;
disk_mem[10726] = 0;
disk_mem[10727] = 0;
disk_mem[10728] = 0;
disk_mem[10729] = 0;
disk_mem[10730] = 0;
disk_mem[10731] = 0;
disk_mem[10732] = 0;
disk_mem[10733] = 0;
disk_mem[10734] = 0;
disk_mem[10735] = 0;
disk_mem[10736] = 0;
disk_mem[10737] = 0;
disk_mem[10738] = 0;
disk_mem[10739] = 0;
disk_mem[10740] = 0;
disk_mem[10741] = 0;
disk_mem[10742] = 0;
disk_mem[10743] = 0;
disk_mem[10744] = 0;
disk_mem[10745] = 0;
disk_mem[10746] = 0;
disk_mem[10747] = 0;
disk_mem[10748] = 0;
disk_mem[10749] = 0;
disk_mem[10750] = 0;
disk_mem[10751] = 0;
disk_mem[10752] = 0;
disk_mem[10753] = 0;
disk_mem[10754] = 0;
disk_mem[10755] = 0;
disk_mem[10756] = 0;
disk_mem[10757] = 0;
disk_mem[10758] = 0;
disk_mem[10759] = 0;
disk_mem[10760] = 0;
disk_mem[10761] = 0;
disk_mem[10762] = 0;
disk_mem[10763] = 0;
disk_mem[10764] = 0;
disk_mem[10765] = 0;
disk_mem[10766] = 0;
disk_mem[10767] = 0;
disk_mem[10768] = 0;
disk_mem[10769] = 0;
disk_mem[10770] = 0;
disk_mem[10771] = 0;
disk_mem[10772] = 0;
disk_mem[10773] = 0;
disk_mem[10774] = 0;
disk_mem[10775] = 0;
disk_mem[10776] = 0;
disk_mem[10777] = 0;
disk_mem[10778] = 0;
disk_mem[10779] = 0;
disk_mem[10780] = 0;
disk_mem[10781] = 0;
disk_mem[10782] = 0;
disk_mem[10783] = 0;
disk_mem[10784] = 0;
disk_mem[10785] = 0;
disk_mem[10786] = 0;
disk_mem[10787] = 0;
disk_mem[10788] = 0;
disk_mem[10789] = 0;
disk_mem[10790] = 0;
disk_mem[10791] = 0;
disk_mem[10792] = 0;
disk_mem[10793] = 0;
disk_mem[10794] = 0;
disk_mem[10795] = 0;
disk_mem[10796] = 0;
disk_mem[10797] = 0;
disk_mem[10798] = 0;
disk_mem[10799] = 0;
disk_mem[10800] = 0;
disk_mem[10801] = 0;
disk_mem[10802] = 0;
disk_mem[10803] = 0;
disk_mem[10804] = 0;
disk_mem[10805] = 0;
disk_mem[10806] = 0;
disk_mem[10807] = 0;
disk_mem[10808] = 0;
disk_mem[10809] = 0;
disk_mem[10810] = 0;
disk_mem[10811] = 0;
disk_mem[10812] = 0;
disk_mem[10813] = 0;
disk_mem[10814] = 0;
disk_mem[10815] = 0;
disk_mem[10816] = 0;
disk_mem[10817] = 0;
disk_mem[10818] = 0;
disk_mem[10819] = 0;
disk_mem[10820] = 0;
disk_mem[10821] = 0;
disk_mem[10822] = 0;
disk_mem[10823] = 0;
disk_mem[10824] = 0;
disk_mem[10825] = 0;
disk_mem[10826] = 0;
disk_mem[10827] = 0;
disk_mem[10828] = 0;
disk_mem[10829] = 0;
disk_mem[10830] = 0;
disk_mem[10831] = 0;
disk_mem[10832] = 0;
disk_mem[10833] = 0;
disk_mem[10834] = 0;
disk_mem[10835] = 0;
disk_mem[10836] = 0;
disk_mem[10837] = 0;
disk_mem[10838] = 0;
disk_mem[10839] = 0;
disk_mem[10840] = 0;
disk_mem[10841] = 0;
disk_mem[10842] = 0;
disk_mem[10843] = 0;
disk_mem[10844] = 0;
disk_mem[10845] = 0;
disk_mem[10846] = 0;
disk_mem[10847] = 0;
disk_mem[10848] = 0;
disk_mem[10849] = 0;
disk_mem[10850] = 0;
disk_mem[10851] = 0;
disk_mem[10852] = 0;
disk_mem[10853] = 0;
disk_mem[10854] = 0;
disk_mem[10855] = 0;
disk_mem[10856] = 0;
disk_mem[10857] = 0;
disk_mem[10858] = 0;
disk_mem[10859] = 0;
disk_mem[10860] = 0;
disk_mem[10861] = 0;
disk_mem[10862] = 0;
disk_mem[10863] = 0;
disk_mem[10864] = 0;
disk_mem[10865] = 0;
disk_mem[10866] = 0;
disk_mem[10867] = 0;
disk_mem[10868] = 0;
disk_mem[10869] = 0;
disk_mem[10870] = 0;
disk_mem[10871] = 0;
disk_mem[10872] = 0;
disk_mem[10873] = 0;
disk_mem[10874] = 0;
disk_mem[10875] = 0;
disk_mem[10876] = 0;
disk_mem[10877] = 0;
disk_mem[10878] = 0;
disk_mem[10879] = 0;
disk_mem[10880] = 0;
disk_mem[10881] = 0;
disk_mem[10882] = 0;
disk_mem[10883] = 0;
disk_mem[10884] = 0;
disk_mem[10885] = 0;
disk_mem[10886] = 0;
disk_mem[10887] = 0;
disk_mem[10888] = 0;
disk_mem[10889] = 0;
disk_mem[10890] = 0;
disk_mem[10891] = 0;
disk_mem[10892] = 0;
disk_mem[10893] = 0;
disk_mem[10894] = 0;
disk_mem[10895] = 0;
disk_mem[10896] = 0;
disk_mem[10897] = 0;
disk_mem[10898] = 0;
disk_mem[10899] = 0;
disk_mem[10900] = 0;
disk_mem[10901] = 0;
disk_mem[10902] = 0;
disk_mem[10903] = 0;
disk_mem[10904] = 0;
disk_mem[10905] = 0;
disk_mem[10906] = 0;
disk_mem[10907] = 0;
disk_mem[10908] = 0;
disk_mem[10909] = 0;
disk_mem[10910] = 0;
disk_mem[10911] = 0;
disk_mem[10912] = 0;
disk_mem[10913] = 0;
disk_mem[10914] = 0;
disk_mem[10915] = 0;
disk_mem[10916] = 0;
disk_mem[10917] = 0;
disk_mem[10918] = 0;
disk_mem[10919] = 0;
disk_mem[10920] = 0;
disk_mem[10921] = 0;
disk_mem[10922] = 0;
disk_mem[10923] = 0;
disk_mem[10924] = 0;
disk_mem[10925] = 0;
disk_mem[10926] = 0;
disk_mem[10927] = 0;
disk_mem[10928] = 0;
disk_mem[10929] = 0;
disk_mem[10930] = 0;
disk_mem[10931] = 0;
disk_mem[10932] = 0;
disk_mem[10933] = 0;
disk_mem[10934] = 0;
disk_mem[10935] = 0;
disk_mem[10936] = 0;
disk_mem[10937] = 0;
disk_mem[10938] = 0;
disk_mem[10939] = 0;
disk_mem[10940] = 0;
disk_mem[10941] = 0;
disk_mem[10942] = 0;
disk_mem[10943] = 0;
disk_mem[10944] = 0;
disk_mem[10945] = 0;
disk_mem[10946] = 0;
disk_mem[10947] = 0;
disk_mem[10948] = 0;
disk_mem[10949] = 0;
disk_mem[10950] = 0;
disk_mem[10951] = 0;
disk_mem[10952] = 0;
disk_mem[10953] = 0;
disk_mem[10954] = 0;
disk_mem[10955] = 0;
disk_mem[10956] = 0;
disk_mem[10957] = 0;
disk_mem[10958] = 0;
disk_mem[10959] = 0;
disk_mem[10960] = 0;
disk_mem[10961] = 0;
disk_mem[10962] = 0;
disk_mem[10963] = 0;
disk_mem[10964] = 0;
disk_mem[10965] = 0;
disk_mem[10966] = 0;
disk_mem[10967] = 0;
disk_mem[10968] = 0;
disk_mem[10969] = 0;
disk_mem[10970] = 0;
disk_mem[10971] = 0;
disk_mem[10972] = 0;
disk_mem[10973] = 0;
disk_mem[10974] = 0;
disk_mem[10975] = 0;
disk_mem[10976] = 0;
disk_mem[10977] = 0;
disk_mem[10978] = 0;
disk_mem[10979] = 0;
disk_mem[10980] = 0;
disk_mem[10981] = 0;
disk_mem[10982] = 0;
disk_mem[10983] = 0;
disk_mem[10984] = 0;
disk_mem[10985] = 0;
disk_mem[10986] = 0;
disk_mem[10987] = 0;
disk_mem[10988] = 0;
disk_mem[10989] = 0;
disk_mem[10990] = 0;
disk_mem[10991] = 0;
disk_mem[10992] = 0;
disk_mem[10993] = 0;
disk_mem[10994] = 0;
disk_mem[10995] = 0;
disk_mem[10996] = 0;
disk_mem[10997] = 0;
disk_mem[10998] = 0;
disk_mem[10999] = 0;
disk_mem[11000] = 0;
disk_mem[11001] = 0;
disk_mem[11002] = 0;
disk_mem[11003] = 0;
disk_mem[11004] = 0;
disk_mem[11005] = 0;
disk_mem[11006] = 0;
disk_mem[11007] = 0;
disk_mem[11008] = 0;
disk_mem[11009] = 0;
disk_mem[11010] = 0;
disk_mem[11011] = 0;
disk_mem[11012] = 0;
disk_mem[11013] = 0;
disk_mem[11014] = 0;
disk_mem[11015] = 0;
disk_mem[11016] = 0;
disk_mem[11017] = 0;
disk_mem[11018] = 0;
disk_mem[11019] = 0;
disk_mem[11020] = 0;
disk_mem[11021] = 0;
disk_mem[11022] = 0;
disk_mem[11023] = 0;
disk_mem[11024] = 0;
disk_mem[11025] = 0;
disk_mem[11026] = 0;
disk_mem[11027] = 0;
disk_mem[11028] = 0;
disk_mem[11029] = 0;
disk_mem[11030] = 0;
disk_mem[11031] = 0;
disk_mem[11032] = 0;
disk_mem[11033] = 0;
disk_mem[11034] = 0;
disk_mem[11035] = 0;
disk_mem[11036] = 0;
disk_mem[11037] = 0;
disk_mem[11038] = 0;
disk_mem[11039] = 0;
disk_mem[11040] = 0;
disk_mem[11041] = 0;
disk_mem[11042] = 0;
disk_mem[11043] = 0;
disk_mem[11044] = 0;
disk_mem[11045] = 0;
disk_mem[11046] = 0;
disk_mem[11047] = 0;
disk_mem[11048] = 0;
disk_mem[11049] = 0;
disk_mem[11050] = 0;
disk_mem[11051] = 0;
disk_mem[11052] = 0;
disk_mem[11053] = 0;
disk_mem[11054] = 0;
disk_mem[11055] = 0;
disk_mem[11056] = 0;
disk_mem[11057] = 0;
disk_mem[11058] = 0;
disk_mem[11059] = 0;
disk_mem[11060] = 0;
disk_mem[11061] = 0;
disk_mem[11062] = 0;
disk_mem[11063] = 0;
disk_mem[11064] = 0;
disk_mem[11065] = 0;
disk_mem[11066] = 0;
disk_mem[11067] = 0;
disk_mem[11068] = 0;
disk_mem[11069] = 0;
disk_mem[11070] = 0;
disk_mem[11071] = 0;
disk_mem[11072] = 0;
disk_mem[11073] = 0;
disk_mem[11074] = 0;
disk_mem[11075] = 0;
disk_mem[11076] = 0;
disk_mem[11077] = 0;
disk_mem[11078] = 0;
disk_mem[11079] = 0;
disk_mem[11080] = 0;
disk_mem[11081] = 0;
disk_mem[11082] = 0;
disk_mem[11083] = 0;
disk_mem[11084] = 0;
disk_mem[11085] = 0;
disk_mem[11086] = 0;
disk_mem[11087] = 0;
disk_mem[11088] = 0;
disk_mem[11089] = 0;
disk_mem[11090] = 0;
disk_mem[11091] = 0;
disk_mem[11092] = 0;
disk_mem[11093] = 0;
disk_mem[11094] = 0;
disk_mem[11095] = 0;
disk_mem[11096] = 0;
disk_mem[11097] = 0;
disk_mem[11098] = 0;
disk_mem[11099] = 0;
disk_mem[11100] = 0;
disk_mem[11101] = 0;
disk_mem[11102] = 0;
disk_mem[11103] = 0;
disk_mem[11104] = 0;
disk_mem[11105] = 0;
disk_mem[11106] = 0;
disk_mem[11107] = 0;
disk_mem[11108] = 0;
disk_mem[11109] = 0;
disk_mem[11110] = 0;
disk_mem[11111] = 0;
disk_mem[11112] = 0;
disk_mem[11113] = 0;
disk_mem[11114] = 0;
disk_mem[11115] = 0;
disk_mem[11116] = 0;
disk_mem[11117] = 0;
disk_mem[11118] = 0;
disk_mem[11119] = 0;
disk_mem[11120] = 0;
disk_mem[11121] = 0;
disk_mem[11122] = 0;
disk_mem[11123] = 0;
disk_mem[11124] = 0;
disk_mem[11125] = 0;
disk_mem[11126] = 0;
disk_mem[11127] = 0;
disk_mem[11128] = 0;
disk_mem[11129] = 0;
disk_mem[11130] = 0;
disk_mem[11131] = 0;
disk_mem[11132] = 0;
disk_mem[11133] = 0;
disk_mem[11134] = 0;
disk_mem[11135] = 0;
disk_mem[11136] = 0;
disk_mem[11137] = 0;
disk_mem[11138] = 0;
disk_mem[11139] = 0;
disk_mem[11140] = 0;
disk_mem[11141] = 0;
disk_mem[11142] = 0;
disk_mem[11143] = 0;
disk_mem[11144] = 0;
disk_mem[11145] = 0;
disk_mem[11146] = 0;
disk_mem[11147] = 0;
disk_mem[11148] = 0;
disk_mem[11149] = 0;
disk_mem[11150] = 0;
disk_mem[11151] = 0;
disk_mem[11152] = 0;
disk_mem[11153] = 0;
disk_mem[11154] = 0;
disk_mem[11155] = 0;
disk_mem[11156] = 0;
disk_mem[11157] = 0;
disk_mem[11158] = 0;
disk_mem[11159] = 0;
disk_mem[11160] = 0;
disk_mem[11161] = 0;
disk_mem[11162] = 0;
disk_mem[11163] = 0;
disk_mem[11164] = 0;
disk_mem[11165] = 0;
disk_mem[11166] = 0;
disk_mem[11167] = 0;
disk_mem[11168] = 0;
disk_mem[11169] = 0;
disk_mem[11170] = 0;
disk_mem[11171] = 0;
disk_mem[11172] = 0;
disk_mem[11173] = 0;
disk_mem[11174] = 0;
disk_mem[11175] = 0;
disk_mem[11176] = 0;
disk_mem[11177] = 0;
disk_mem[11178] = 0;
disk_mem[11179] = 0;
disk_mem[11180] = 0;
disk_mem[11181] = 0;
disk_mem[11182] = 0;
disk_mem[11183] = 0;
disk_mem[11184] = 0;
disk_mem[11185] = 0;
disk_mem[11186] = 0;
disk_mem[11187] = 0;
disk_mem[11188] = 0;
disk_mem[11189] = 0;
disk_mem[11190] = 0;
disk_mem[11191] = 0;
disk_mem[11192] = 0;
disk_mem[11193] = 0;
disk_mem[11194] = 0;
disk_mem[11195] = 0;
disk_mem[11196] = 0;
disk_mem[11197] = 0;
disk_mem[11198] = 0;
disk_mem[11199] = 0;
disk_mem[11200] = 0;
disk_mem[11201] = 0;
disk_mem[11202] = 0;
disk_mem[11203] = 0;
disk_mem[11204] = 0;
disk_mem[11205] = 0;
disk_mem[11206] = 0;
disk_mem[11207] = 0;
disk_mem[11208] = 0;
disk_mem[11209] = 0;
disk_mem[11210] = 0;
disk_mem[11211] = 0;
disk_mem[11212] = 0;
disk_mem[11213] = 0;
disk_mem[11214] = 0;
disk_mem[11215] = 0;
disk_mem[11216] = 0;
disk_mem[11217] = 0;
disk_mem[11218] = 0;
disk_mem[11219] = 0;
disk_mem[11220] = 0;
disk_mem[11221] = 0;
disk_mem[11222] = 0;
disk_mem[11223] = 0;
disk_mem[11224] = 0;
disk_mem[11225] = 0;
disk_mem[11226] = 0;
disk_mem[11227] = 0;
disk_mem[11228] = 0;
disk_mem[11229] = 0;
disk_mem[11230] = 0;
disk_mem[11231] = 0;
disk_mem[11232] = 0;
disk_mem[11233] = 0;
disk_mem[11234] = 0;
disk_mem[11235] = 0;
disk_mem[11236] = 0;
disk_mem[11237] = 0;
disk_mem[11238] = 0;
disk_mem[11239] = 0;
disk_mem[11240] = 0;
disk_mem[11241] = 0;
disk_mem[11242] = 0;
disk_mem[11243] = 0;
disk_mem[11244] = 0;
disk_mem[11245] = 0;
disk_mem[11246] = 0;
disk_mem[11247] = 0;
disk_mem[11248] = 0;
disk_mem[11249] = 0;
disk_mem[11250] = 0;
disk_mem[11251] = 0;
disk_mem[11252] = 0;
disk_mem[11253] = 0;
disk_mem[11254] = 0;
disk_mem[11255] = 0;
disk_mem[11256] = 0;
disk_mem[11257] = 0;
disk_mem[11258] = 0;
disk_mem[11259] = 0;
disk_mem[11260] = 0;
disk_mem[11261] = 0;
disk_mem[11262] = 0;
disk_mem[11263] = 0;
disk_mem[11264] = 0;
disk_mem[11265] = 0;
disk_mem[11266] = 0;
disk_mem[11267] = 0;
disk_mem[11268] = 0;
disk_mem[11269] = 0;
disk_mem[11270] = 0;
disk_mem[11271] = 0;
disk_mem[11272] = 0;
disk_mem[11273] = 0;
disk_mem[11274] = 0;
disk_mem[11275] = 0;
disk_mem[11276] = 0;
disk_mem[11277] = 0;
disk_mem[11278] = 0;
disk_mem[11279] = 0;
disk_mem[11280] = 0;
disk_mem[11281] = 0;
disk_mem[11282] = 0;
disk_mem[11283] = 0;
disk_mem[11284] = 0;
disk_mem[11285] = 0;
disk_mem[11286] = 0;
disk_mem[11287] = 0;
disk_mem[11288] = 0;
disk_mem[11289] = 0;
disk_mem[11290] = 0;
disk_mem[11291] = 0;
disk_mem[11292] = 0;
disk_mem[11293] = 0;
disk_mem[11294] = 0;
disk_mem[11295] = 0;
disk_mem[11296] = 0;
disk_mem[11297] = 0;
disk_mem[11298] = 0;
disk_mem[11299] = 0;
disk_mem[11300] = 0;
disk_mem[11301] = 0;
disk_mem[11302] = 0;
disk_mem[11303] = 0;
disk_mem[11304] = 0;
disk_mem[11305] = 0;
disk_mem[11306] = 0;
disk_mem[11307] = 0;
disk_mem[11308] = 0;
disk_mem[11309] = 0;
disk_mem[11310] = 0;
disk_mem[11311] = 0;
disk_mem[11312] = 0;
disk_mem[11313] = 0;
disk_mem[11314] = 0;
disk_mem[11315] = 0;
disk_mem[11316] = 0;
disk_mem[11317] = 0;
disk_mem[11318] = 0;
disk_mem[11319] = 0;
disk_mem[11320] = 0;
disk_mem[11321] = 0;
disk_mem[11322] = 0;
disk_mem[11323] = 0;
disk_mem[11324] = 0;
disk_mem[11325] = 0;
disk_mem[11326] = 0;
disk_mem[11327] = 0;
disk_mem[11328] = 0;
disk_mem[11329] = 0;
disk_mem[11330] = 0;
disk_mem[11331] = 0;
disk_mem[11332] = 0;
disk_mem[11333] = 0;
disk_mem[11334] = 0;
disk_mem[11335] = 0;
disk_mem[11336] = 0;
disk_mem[11337] = 0;
disk_mem[11338] = 0;
disk_mem[11339] = 0;
disk_mem[11340] = 0;
disk_mem[11341] = 0;
disk_mem[11342] = 0;
disk_mem[11343] = 0;
disk_mem[11344] = 0;
disk_mem[11345] = 0;
disk_mem[11346] = 0;
disk_mem[11347] = 0;
disk_mem[11348] = 0;
disk_mem[11349] = 0;
disk_mem[11350] = 0;
disk_mem[11351] = 0;
disk_mem[11352] = 0;
disk_mem[11353] = 0;
disk_mem[11354] = 0;
disk_mem[11355] = 0;
disk_mem[11356] = 0;
disk_mem[11357] = 0;
disk_mem[11358] = 0;
disk_mem[11359] = 0;
disk_mem[11360] = 0;
disk_mem[11361] = 0;
disk_mem[11362] = 0;
disk_mem[11363] = 0;
disk_mem[11364] = 0;
disk_mem[11365] = 0;
disk_mem[11366] = 0;
disk_mem[11367] = 0;
disk_mem[11368] = 0;
disk_mem[11369] = 0;
disk_mem[11370] = 0;
disk_mem[11371] = 0;
disk_mem[11372] = 0;
disk_mem[11373] = 0;
disk_mem[11374] = 0;
disk_mem[11375] = 0;
disk_mem[11376] = 0;
disk_mem[11377] = 0;
disk_mem[11378] = 0;
disk_mem[11379] = 0;
disk_mem[11380] = 0;
disk_mem[11381] = 0;
disk_mem[11382] = 0;
disk_mem[11383] = 0;
disk_mem[11384] = 0;
disk_mem[11385] = 0;
disk_mem[11386] = 0;
disk_mem[11387] = 0;
disk_mem[11388] = 0;
disk_mem[11389] = 0;
disk_mem[11390] = 0;
disk_mem[11391] = 0;
disk_mem[11392] = 0;
disk_mem[11393] = 0;
disk_mem[11394] = 0;
disk_mem[11395] = 0;
disk_mem[11396] = 0;
disk_mem[11397] = 0;
disk_mem[11398] = 0;
disk_mem[11399] = 0;
disk_mem[11400] = 0;
disk_mem[11401] = 0;
disk_mem[11402] = 0;
disk_mem[11403] = 0;
disk_mem[11404] = 0;
disk_mem[11405] = 0;
disk_mem[11406] = 0;
disk_mem[11407] = 0;
disk_mem[11408] = 0;
disk_mem[11409] = 0;
disk_mem[11410] = 0;
disk_mem[11411] = 0;
disk_mem[11412] = 0;
disk_mem[11413] = 0;
disk_mem[11414] = 0;
disk_mem[11415] = 0;
disk_mem[11416] = 0;
disk_mem[11417] = 0;
disk_mem[11418] = 0;
disk_mem[11419] = 0;
disk_mem[11420] = 0;
disk_mem[11421] = 0;
disk_mem[11422] = 0;
disk_mem[11423] = 0;
disk_mem[11424] = 0;
disk_mem[11425] = 0;
disk_mem[11426] = 0;
disk_mem[11427] = 0;
disk_mem[11428] = 0;
disk_mem[11429] = 0;
disk_mem[11430] = 0;
disk_mem[11431] = 0;
disk_mem[11432] = 0;
disk_mem[11433] = 0;
disk_mem[11434] = 0;
disk_mem[11435] = 0;
disk_mem[11436] = 0;
disk_mem[11437] = 0;
disk_mem[11438] = 0;
disk_mem[11439] = 0;
disk_mem[11440] = 0;
disk_mem[11441] = 0;
disk_mem[11442] = 0;
disk_mem[11443] = 0;
disk_mem[11444] = 0;
disk_mem[11445] = 0;
disk_mem[11446] = 0;
disk_mem[11447] = 0;
disk_mem[11448] = 0;
disk_mem[11449] = 0;
disk_mem[11450] = 0;
disk_mem[11451] = 0;
disk_mem[11452] = 0;
disk_mem[11453] = 0;
disk_mem[11454] = 0;
disk_mem[11455] = 0;
disk_mem[11456] = 0;
disk_mem[11457] = 0;
disk_mem[11458] = 0;
disk_mem[11459] = 0;
disk_mem[11460] = 0;
disk_mem[11461] = 0;
disk_mem[11462] = 0;
disk_mem[11463] = 0;
disk_mem[11464] = 0;
disk_mem[11465] = 0;
disk_mem[11466] = 0;
disk_mem[11467] = 0;
disk_mem[11468] = 0;
disk_mem[11469] = 0;
disk_mem[11470] = 0;
disk_mem[11471] = 0;
disk_mem[11472] = 0;
disk_mem[11473] = 0;
disk_mem[11474] = 0;
disk_mem[11475] = 0;
disk_mem[11476] = 0;
disk_mem[11477] = 0;
disk_mem[11478] = 0;
disk_mem[11479] = 0;
disk_mem[11480] = 0;
disk_mem[11481] = 0;
disk_mem[11482] = 0;
disk_mem[11483] = 0;
disk_mem[11484] = 0;
disk_mem[11485] = 0;
disk_mem[11486] = 0;
disk_mem[11487] = 0;
disk_mem[11488] = 0;
disk_mem[11489] = 0;
disk_mem[11490] = 0;
disk_mem[11491] = 0;
disk_mem[11492] = 0;
disk_mem[11493] = 0;
disk_mem[11494] = 0;
disk_mem[11495] = 0;
disk_mem[11496] = 0;
disk_mem[11497] = 0;
disk_mem[11498] = 0;
disk_mem[11499] = 0;
disk_mem[11500] = 0;
disk_mem[11501] = 0;
disk_mem[11502] = 0;
disk_mem[11503] = 0;
disk_mem[11504] = 0;
disk_mem[11505] = 0;
disk_mem[11506] = 0;
disk_mem[11507] = 0;
disk_mem[11508] = 0;
disk_mem[11509] = 0;
disk_mem[11510] = 0;
disk_mem[11511] = 0;
disk_mem[11512] = 0;
disk_mem[11513] = 0;
disk_mem[11514] = 0;
disk_mem[11515] = 0;
disk_mem[11516] = 0;
disk_mem[11517] = 0;
disk_mem[11518] = 0;
disk_mem[11519] = 0;
disk_mem[11520] = 0;
disk_mem[11521] = 0;
disk_mem[11522] = 0;
disk_mem[11523] = 0;
disk_mem[11524] = 0;
disk_mem[11525] = 0;
disk_mem[11526] = 0;
disk_mem[11527] = 0;
disk_mem[11528] = 0;
disk_mem[11529] = 0;
disk_mem[11530] = 0;
disk_mem[11531] = 0;
disk_mem[11532] = 0;
disk_mem[11533] = 0;
disk_mem[11534] = 0;
disk_mem[11535] = 0;
disk_mem[11536] = 0;
disk_mem[11537] = 0;
disk_mem[11538] = 0;
disk_mem[11539] = 0;
disk_mem[11540] = 0;
disk_mem[11541] = 0;
disk_mem[11542] = 0;
disk_mem[11543] = 0;
disk_mem[11544] = 0;
disk_mem[11545] = 0;
disk_mem[11546] = 0;
disk_mem[11547] = 0;
disk_mem[11548] = 0;
disk_mem[11549] = 0;
disk_mem[11550] = 0;
disk_mem[11551] = 0;
disk_mem[11552] = 0;
disk_mem[11553] = 0;
disk_mem[11554] = 0;
disk_mem[11555] = 0;
disk_mem[11556] = 0;
disk_mem[11557] = 0;
disk_mem[11558] = 0;
disk_mem[11559] = 0;
disk_mem[11560] = 0;
disk_mem[11561] = 0;
disk_mem[11562] = 0;
disk_mem[11563] = 0;
disk_mem[11564] = 0;
disk_mem[11565] = 0;
disk_mem[11566] = 0;
disk_mem[11567] = 0;
disk_mem[11568] = 0;
disk_mem[11569] = 0;
disk_mem[11570] = 0;
disk_mem[11571] = 0;
disk_mem[11572] = 0;
disk_mem[11573] = 0;
disk_mem[11574] = 0;
disk_mem[11575] = 0;
disk_mem[11576] = 0;
disk_mem[11577] = 0;
disk_mem[11578] = 0;
disk_mem[11579] = 0;
disk_mem[11580] = 0;
disk_mem[11581] = 0;
disk_mem[11582] = 0;
disk_mem[11583] = 0;
disk_mem[11584] = 0;
disk_mem[11585] = 0;
disk_mem[11586] = 0;
disk_mem[11587] = 0;
disk_mem[11588] = 0;
disk_mem[11589] = 0;
disk_mem[11590] = 0;
disk_mem[11591] = 0;
disk_mem[11592] = 0;
disk_mem[11593] = 0;
disk_mem[11594] = 0;
disk_mem[11595] = 0;
disk_mem[11596] = 0;
disk_mem[11597] = 0;
disk_mem[11598] = 0;
disk_mem[11599] = 0;
disk_mem[11600] = 0;
disk_mem[11601] = 0;
disk_mem[11602] = 0;
disk_mem[11603] = 0;
disk_mem[11604] = 0;
disk_mem[11605] = 0;
disk_mem[11606] = 0;
disk_mem[11607] = 0;
disk_mem[11608] = 0;
disk_mem[11609] = 0;
disk_mem[11610] = 0;
disk_mem[11611] = 0;
disk_mem[11612] = 0;
disk_mem[11613] = 0;
disk_mem[11614] = 0;
disk_mem[11615] = 0;
disk_mem[11616] = 0;
disk_mem[11617] = 0;
disk_mem[11618] = 0;
disk_mem[11619] = 0;
disk_mem[11620] = 0;
disk_mem[11621] = 0;
disk_mem[11622] = 0;
disk_mem[11623] = 0;
disk_mem[11624] = 0;
disk_mem[11625] = 0;
disk_mem[11626] = 0;
disk_mem[11627] = 0;
disk_mem[11628] = 0;
disk_mem[11629] = 0;
disk_mem[11630] = 0;
disk_mem[11631] = 0;
disk_mem[11632] = 0;
disk_mem[11633] = 0;
disk_mem[11634] = 0;
disk_mem[11635] = 0;
disk_mem[11636] = 0;
disk_mem[11637] = 0;
disk_mem[11638] = 0;
disk_mem[11639] = 0;
disk_mem[11640] = 0;
disk_mem[11641] = 0;
disk_mem[11642] = 0;
disk_mem[11643] = 0;
disk_mem[11644] = 0;
disk_mem[11645] = 0;
disk_mem[11646] = 0;
disk_mem[11647] = 0;
disk_mem[11648] = 0;
disk_mem[11649] = 0;
disk_mem[11650] = 0;
disk_mem[11651] = 0;
disk_mem[11652] = 0;
disk_mem[11653] = 0;
disk_mem[11654] = 0;
disk_mem[11655] = 0;
disk_mem[11656] = 0;
disk_mem[11657] = 0;
disk_mem[11658] = 0;
disk_mem[11659] = 0;
disk_mem[11660] = 0;
disk_mem[11661] = 0;
disk_mem[11662] = 0;
disk_mem[11663] = 0;
disk_mem[11664] = 0;
disk_mem[11665] = 0;
disk_mem[11666] = 0;
disk_mem[11667] = 0;
disk_mem[11668] = 0;
disk_mem[11669] = 0;
disk_mem[11670] = 0;
disk_mem[11671] = 0;
disk_mem[11672] = 0;
disk_mem[11673] = 0;
disk_mem[11674] = 0;
disk_mem[11675] = 0;
disk_mem[11676] = 0;
disk_mem[11677] = 0;
disk_mem[11678] = 0;
disk_mem[11679] = 0;
disk_mem[11680] = 0;
disk_mem[11681] = 0;
disk_mem[11682] = 0;
disk_mem[11683] = 0;
disk_mem[11684] = 0;
disk_mem[11685] = 0;
disk_mem[11686] = 0;
disk_mem[11687] = 0;
disk_mem[11688] = 0;
disk_mem[11689] = 0;
disk_mem[11690] = 0;
disk_mem[11691] = 0;
disk_mem[11692] = 0;
disk_mem[11693] = 0;
disk_mem[11694] = 0;
disk_mem[11695] = 0;
disk_mem[11696] = 0;
disk_mem[11697] = 0;
disk_mem[11698] = 0;
disk_mem[11699] = 0;
disk_mem[11700] = 0;
disk_mem[11701] = 0;
disk_mem[11702] = 0;
disk_mem[11703] = 0;
disk_mem[11704] = 0;
disk_mem[11705] = 0;
disk_mem[11706] = 0;
disk_mem[11707] = 0;
disk_mem[11708] = 0;
disk_mem[11709] = 0;
disk_mem[11710] = 0;
disk_mem[11711] = 0;
disk_mem[11712] = 0;
disk_mem[11713] = 0;
disk_mem[11714] = 0;
disk_mem[11715] = 0;
disk_mem[11716] = 0;
disk_mem[11717] = 0;
disk_mem[11718] = 0;
disk_mem[11719] = 0;
disk_mem[11720] = 0;
disk_mem[11721] = 0;
disk_mem[11722] = 0;
disk_mem[11723] = 0;
disk_mem[11724] = 0;
disk_mem[11725] = 0;
disk_mem[11726] = 0;
disk_mem[11727] = 0;
disk_mem[11728] = 0;
disk_mem[11729] = 0;
disk_mem[11730] = 0;
disk_mem[11731] = 0;
disk_mem[11732] = 0;
disk_mem[11733] = 0;
disk_mem[11734] = 0;
disk_mem[11735] = 0;
disk_mem[11736] = 0;
disk_mem[11737] = 0;
disk_mem[11738] = 0;
disk_mem[11739] = 0;
disk_mem[11740] = 0;
disk_mem[11741] = 0;
disk_mem[11742] = 0;
disk_mem[11743] = 0;
disk_mem[11744] = 0;
disk_mem[11745] = 0;
disk_mem[11746] = 0;
disk_mem[11747] = 0;
disk_mem[11748] = 0;
disk_mem[11749] = 0;
disk_mem[11750] = 0;
disk_mem[11751] = 0;
disk_mem[11752] = 0;
disk_mem[11753] = 0;
disk_mem[11754] = 0;
disk_mem[11755] = 0;
disk_mem[11756] = 0;
disk_mem[11757] = 0;
disk_mem[11758] = 0;
disk_mem[11759] = 0;
disk_mem[11760] = 0;
disk_mem[11761] = 0;
disk_mem[11762] = 0;
disk_mem[11763] = 0;
disk_mem[11764] = 0;
disk_mem[11765] = 0;
disk_mem[11766] = 0;
disk_mem[11767] = 0;
disk_mem[11768] = 0;
disk_mem[11769] = 0;
disk_mem[11770] = 0;
disk_mem[11771] = 0;
disk_mem[11772] = 0;
disk_mem[11773] = 0;
disk_mem[11774] = 0;
disk_mem[11775] = 0;
disk_mem[11776] = 0;
disk_mem[11777] = 0;
disk_mem[11778] = 0;
disk_mem[11779] = 0;
disk_mem[11780] = 0;
disk_mem[11781] = 0;
disk_mem[11782] = 0;
disk_mem[11783] = 0;
disk_mem[11784] = 0;
disk_mem[11785] = 0;
disk_mem[11786] = 0;
disk_mem[11787] = 0;
disk_mem[11788] = 0;
disk_mem[11789] = 0;
disk_mem[11790] = 0;
disk_mem[11791] = 0;
disk_mem[11792] = 0;
disk_mem[11793] = 0;
disk_mem[11794] = 0;
disk_mem[11795] = 0;
disk_mem[11796] = 0;
disk_mem[11797] = 0;
disk_mem[11798] = 0;
disk_mem[11799] = 0;
disk_mem[11800] = 0;
disk_mem[11801] = 0;
disk_mem[11802] = 0;
disk_mem[11803] = 0;
disk_mem[11804] = 0;
disk_mem[11805] = 0;
disk_mem[11806] = 0;
disk_mem[11807] = 0;
disk_mem[11808] = 0;
disk_mem[11809] = 0;
disk_mem[11810] = 0;
disk_mem[11811] = 0;
disk_mem[11812] = 0;
disk_mem[11813] = 0;
disk_mem[11814] = 0;
disk_mem[11815] = 0;
disk_mem[11816] = 0;
disk_mem[11817] = 0;
disk_mem[11818] = 0;
disk_mem[11819] = 0;
disk_mem[11820] = 0;
disk_mem[11821] = 0;
disk_mem[11822] = 0;
disk_mem[11823] = 0;
disk_mem[11824] = 0;
disk_mem[11825] = 0;
disk_mem[11826] = 0;
disk_mem[11827] = 0;
disk_mem[11828] = 0;
disk_mem[11829] = 0;
disk_mem[11830] = 0;
disk_mem[11831] = 0;
disk_mem[11832] = 0;
disk_mem[11833] = 0;
disk_mem[11834] = 0;
disk_mem[11835] = 0;
disk_mem[11836] = 0;
disk_mem[11837] = 0;
disk_mem[11838] = 0;
disk_mem[11839] = 0;
disk_mem[11840] = 0;
disk_mem[11841] = 0;
disk_mem[11842] = 0;
disk_mem[11843] = 0;
disk_mem[11844] = 0;
disk_mem[11845] = 0;
disk_mem[11846] = 0;
disk_mem[11847] = 0;
disk_mem[11848] = 0;
disk_mem[11849] = 0;
disk_mem[11850] = 0;
disk_mem[11851] = 0;
disk_mem[11852] = 0;
disk_mem[11853] = 0;
disk_mem[11854] = 0;
disk_mem[11855] = 0;
disk_mem[11856] = 0;
disk_mem[11857] = 0;
disk_mem[11858] = 0;
disk_mem[11859] = 0;
disk_mem[11860] = 0;
disk_mem[11861] = 0;
disk_mem[11862] = 0;
disk_mem[11863] = 0;
disk_mem[11864] = 0;
disk_mem[11865] = 0;
disk_mem[11866] = 0;
disk_mem[11867] = 0;
disk_mem[11868] = 0;
disk_mem[11869] = 0;
disk_mem[11870] = 0;
disk_mem[11871] = 0;
disk_mem[11872] = 0;
disk_mem[11873] = 0;
disk_mem[11874] = 0;
disk_mem[11875] = 0;
disk_mem[11876] = 0;
disk_mem[11877] = 0;
disk_mem[11878] = 0;
disk_mem[11879] = 0;
disk_mem[11880] = 0;
disk_mem[11881] = 0;
disk_mem[11882] = 0;
disk_mem[11883] = 0;
disk_mem[11884] = 0;
disk_mem[11885] = 0;
disk_mem[11886] = 0;
disk_mem[11887] = 0;
disk_mem[11888] = 0;
disk_mem[11889] = 0;
disk_mem[11890] = 0;
disk_mem[11891] = 0;
disk_mem[11892] = 0;
disk_mem[11893] = 0;
disk_mem[11894] = 0;
disk_mem[11895] = 0;
disk_mem[11896] = 0;
disk_mem[11897] = 0;
disk_mem[11898] = 0;
disk_mem[11899] = 0;
disk_mem[11900] = 0;
disk_mem[11901] = 0;
disk_mem[11902] = 0;
disk_mem[11903] = 0;
disk_mem[11904] = 0;
disk_mem[11905] = 0;
disk_mem[11906] = 0;
disk_mem[11907] = 0;
disk_mem[11908] = 0;
disk_mem[11909] = 0;
disk_mem[11910] = 0;
disk_mem[11911] = 0;
disk_mem[11912] = 0;
disk_mem[11913] = 0;
disk_mem[11914] = 0;
disk_mem[11915] = 0;
disk_mem[11916] = 0;
disk_mem[11917] = 0;
disk_mem[11918] = 0;
disk_mem[11919] = 0;
disk_mem[11920] = 0;
disk_mem[11921] = 0;
disk_mem[11922] = 0;
disk_mem[11923] = 0;
disk_mem[11924] = 0;
disk_mem[11925] = 0;
disk_mem[11926] = 0;
disk_mem[11927] = 0;
disk_mem[11928] = 0;
disk_mem[11929] = 0;
disk_mem[11930] = 0;
disk_mem[11931] = 0;
disk_mem[11932] = 0;
disk_mem[11933] = 0;
disk_mem[11934] = 0;
disk_mem[11935] = 0;
disk_mem[11936] = 0;
disk_mem[11937] = 0;
disk_mem[11938] = 0;
disk_mem[11939] = 0;
disk_mem[11940] = 0;
disk_mem[11941] = 0;
disk_mem[11942] = 0;
disk_mem[11943] = 0;
disk_mem[11944] = 0;
disk_mem[11945] = 0;
disk_mem[11946] = 0;
disk_mem[11947] = 0;
disk_mem[11948] = 0;
disk_mem[11949] = 0;
disk_mem[11950] = 0;
disk_mem[11951] = 0;
disk_mem[11952] = 0;
disk_mem[11953] = 0;
disk_mem[11954] = 0;
disk_mem[11955] = 0;
disk_mem[11956] = 0;
disk_mem[11957] = 0;
disk_mem[11958] = 0;
disk_mem[11959] = 0;
disk_mem[11960] = 0;
disk_mem[11961] = 0;
disk_mem[11962] = 0;
disk_mem[11963] = 0;
disk_mem[11964] = 0;
disk_mem[11965] = 0;
disk_mem[11966] = 0;
disk_mem[11967] = 0;
disk_mem[11968] = 0;
disk_mem[11969] = 0;
disk_mem[11970] = 0;
disk_mem[11971] = 0;
disk_mem[11972] = 0;
disk_mem[11973] = 0;
disk_mem[11974] = 0;
disk_mem[11975] = 0;
disk_mem[11976] = 0;
disk_mem[11977] = 0;
disk_mem[11978] = 0;
disk_mem[11979] = 0;
disk_mem[11980] = 0;
disk_mem[11981] = 0;
disk_mem[11982] = 0;
disk_mem[11983] = 0;
disk_mem[11984] = 0;
disk_mem[11985] = 0;
disk_mem[11986] = 0;
disk_mem[11987] = 0;
disk_mem[11988] = 0;
disk_mem[11989] = 0;
disk_mem[11990] = 0;
disk_mem[11991] = 0;
disk_mem[11992] = 0;
disk_mem[11993] = 0;
disk_mem[11994] = 0;
disk_mem[11995] = 0;
disk_mem[11996] = 0;
disk_mem[11997] = 0;
disk_mem[11998] = 0;
disk_mem[11999] = 0;
disk_mem[12000] = 0;
disk_mem[12001] = 0;
disk_mem[12002] = 0;
disk_mem[12003] = 0;
disk_mem[12004] = 0;
disk_mem[12005] = 0;
disk_mem[12006] = 0;
disk_mem[12007] = 0;
disk_mem[12008] = 0;
disk_mem[12009] = 0;
disk_mem[12010] = 0;
disk_mem[12011] = 0;
disk_mem[12012] = 0;
disk_mem[12013] = 0;
disk_mem[12014] = 0;
disk_mem[12015] = 0;
disk_mem[12016] = 0;
disk_mem[12017] = 0;
disk_mem[12018] = 0;
disk_mem[12019] = 0;
disk_mem[12020] = 0;
disk_mem[12021] = 0;
disk_mem[12022] = 0;
disk_mem[12023] = 0;
disk_mem[12024] = 0;
disk_mem[12025] = 0;
disk_mem[12026] = 0;
disk_mem[12027] = 0;
disk_mem[12028] = 0;
disk_mem[12029] = 0;
disk_mem[12030] = 0;
disk_mem[12031] = 0;
disk_mem[12032] = 0;
disk_mem[12033] = 0;
disk_mem[12034] = 0;
disk_mem[12035] = 0;
disk_mem[12036] = 0;
disk_mem[12037] = 0;
disk_mem[12038] = 0;
disk_mem[12039] = 0;
disk_mem[12040] = 0;
disk_mem[12041] = 0;
disk_mem[12042] = 0;
disk_mem[12043] = 0;
disk_mem[12044] = 0;
disk_mem[12045] = 0;
disk_mem[12046] = 0;
disk_mem[12047] = 0;
disk_mem[12048] = 0;
disk_mem[12049] = 0;
disk_mem[12050] = 0;
disk_mem[12051] = 0;
disk_mem[12052] = 0;
disk_mem[12053] = 0;
disk_mem[12054] = 0;
disk_mem[12055] = 0;
disk_mem[12056] = 0;
disk_mem[12057] = 0;
disk_mem[12058] = 0;
disk_mem[12059] = 0;
disk_mem[12060] = 0;
disk_mem[12061] = 0;
disk_mem[12062] = 0;
disk_mem[12063] = 0;
disk_mem[12064] = 0;
disk_mem[12065] = 0;
disk_mem[12066] = 0;
disk_mem[12067] = 0;
disk_mem[12068] = 0;
disk_mem[12069] = 0;
disk_mem[12070] = 0;
disk_mem[12071] = 0;
disk_mem[12072] = 0;
disk_mem[12073] = 0;
disk_mem[12074] = 0;
disk_mem[12075] = 0;
disk_mem[12076] = 0;
disk_mem[12077] = 0;
disk_mem[12078] = 0;
disk_mem[12079] = 0;
disk_mem[12080] = 0;
disk_mem[12081] = 0;
disk_mem[12082] = 0;
disk_mem[12083] = 0;
disk_mem[12084] = 0;
disk_mem[12085] = 0;
disk_mem[12086] = 0;
disk_mem[12087] = 0;
disk_mem[12088] = 0;
disk_mem[12089] = 0;
disk_mem[12090] = 0;
disk_mem[12091] = 0;
disk_mem[12092] = 0;
disk_mem[12093] = 0;
disk_mem[12094] = 0;
disk_mem[12095] = 0;
disk_mem[12096] = 0;
disk_mem[12097] = 0;
disk_mem[12098] = 0;
disk_mem[12099] = 0;
disk_mem[12100] = 0;
disk_mem[12101] = 0;
disk_mem[12102] = 0;
disk_mem[12103] = 0;
disk_mem[12104] = 0;
disk_mem[12105] = 0;
disk_mem[12106] = 0;
disk_mem[12107] = 0;
disk_mem[12108] = 0;
disk_mem[12109] = 0;
disk_mem[12110] = 0;
disk_mem[12111] = 0;
disk_mem[12112] = 0;
disk_mem[12113] = 0;
disk_mem[12114] = 0;
disk_mem[12115] = 0;
disk_mem[12116] = 0;
disk_mem[12117] = 0;
disk_mem[12118] = 0;
disk_mem[12119] = 0;
disk_mem[12120] = 0;
disk_mem[12121] = 0;
disk_mem[12122] = 0;
disk_mem[12123] = 0;
disk_mem[12124] = 0;
disk_mem[12125] = 0;
disk_mem[12126] = 0;
disk_mem[12127] = 0;
disk_mem[12128] = 0;
disk_mem[12129] = 0;
disk_mem[12130] = 0;
disk_mem[12131] = 0;
disk_mem[12132] = 0;
disk_mem[12133] = 0;
disk_mem[12134] = 0;
disk_mem[12135] = 0;
disk_mem[12136] = 0;
disk_mem[12137] = 0;
disk_mem[12138] = 0;
disk_mem[12139] = 0;
disk_mem[12140] = 0;
disk_mem[12141] = 0;
disk_mem[12142] = 0;
disk_mem[12143] = 0;
disk_mem[12144] = 0;
disk_mem[12145] = 0;
disk_mem[12146] = 0;
disk_mem[12147] = 0;
disk_mem[12148] = 0;
disk_mem[12149] = 0;
disk_mem[12150] = 0;
disk_mem[12151] = 0;
disk_mem[12152] = 0;
disk_mem[12153] = 0;
disk_mem[12154] = 0;
disk_mem[12155] = 0;
disk_mem[12156] = 0;
disk_mem[12157] = 0;
disk_mem[12158] = 0;
disk_mem[12159] = 0;
disk_mem[12160] = 0;
disk_mem[12161] = 0;
disk_mem[12162] = 0;
disk_mem[12163] = 0;
disk_mem[12164] = 0;
disk_mem[12165] = 0;
disk_mem[12166] = 0;
disk_mem[12167] = 0;
disk_mem[12168] = 0;
disk_mem[12169] = 0;
disk_mem[12170] = 0;
disk_mem[12171] = 0;
disk_mem[12172] = 0;
disk_mem[12173] = 0;
disk_mem[12174] = 0;
disk_mem[12175] = 0;
disk_mem[12176] = 0;
disk_mem[12177] = 0;
disk_mem[12178] = 0;
disk_mem[12179] = 0;
disk_mem[12180] = 0;
disk_mem[12181] = 0;
disk_mem[12182] = 0;
disk_mem[12183] = 0;
disk_mem[12184] = 0;
disk_mem[12185] = 0;
disk_mem[12186] = 0;
disk_mem[12187] = 0;
disk_mem[12188] = 0;
disk_mem[12189] = 0;
disk_mem[12190] = 0;
disk_mem[12191] = 0;
disk_mem[12192] = 0;
disk_mem[12193] = 0;
disk_mem[12194] = 0;
disk_mem[12195] = 0;
disk_mem[12196] = 0;
disk_mem[12197] = 0;
disk_mem[12198] = 0;
disk_mem[12199] = 0;
disk_mem[12200] = 0;
disk_mem[12201] = 0;
disk_mem[12202] = 0;
disk_mem[12203] = 0;
disk_mem[12204] = 0;
disk_mem[12205] = 0;
disk_mem[12206] = 0;
disk_mem[12207] = 0;
disk_mem[12208] = 0;
disk_mem[12209] = 0;
disk_mem[12210] = 0;
disk_mem[12211] = 0;
disk_mem[12212] = 0;
disk_mem[12213] = 0;
disk_mem[12214] = 0;
disk_mem[12215] = 0;
disk_mem[12216] = 0;
disk_mem[12217] = 0;
disk_mem[12218] = 0;
disk_mem[12219] = 0;
disk_mem[12220] = 0;
disk_mem[12221] = 0;
disk_mem[12222] = 0;
disk_mem[12223] = 0;
disk_mem[12224] = 0;
disk_mem[12225] = 0;
disk_mem[12226] = 0;
disk_mem[12227] = 0;
disk_mem[12228] = 0;
disk_mem[12229] = 0;
disk_mem[12230] = 0;
disk_mem[12231] = 0;
disk_mem[12232] = 0;
disk_mem[12233] = 0;
disk_mem[12234] = 0;
disk_mem[12235] = 0;
disk_mem[12236] = 0;
disk_mem[12237] = 0;
disk_mem[12238] = 0;
disk_mem[12239] = 0;
disk_mem[12240] = 0;
disk_mem[12241] = 0;
disk_mem[12242] = 0;
disk_mem[12243] = 0;
disk_mem[12244] = 0;
disk_mem[12245] = 0;
disk_mem[12246] = 0;
disk_mem[12247] = 0;
disk_mem[12248] = 0;
disk_mem[12249] = 0;
disk_mem[12250] = 0;
disk_mem[12251] = 0;
disk_mem[12252] = 0;
disk_mem[12253] = 0;
disk_mem[12254] = 0;
disk_mem[12255] = 0;
disk_mem[12256] = 0;
disk_mem[12257] = 0;
disk_mem[12258] = 0;
disk_mem[12259] = 0;
disk_mem[12260] = 0;
disk_mem[12261] = 0;
disk_mem[12262] = 0;
disk_mem[12263] = 0;
disk_mem[12264] = 0;
disk_mem[12265] = 0;
disk_mem[12266] = 0;
disk_mem[12267] = 0;
disk_mem[12268] = 0;
disk_mem[12269] = 0;
disk_mem[12270] = 0;
disk_mem[12271] = 0;
disk_mem[12272] = 0;
disk_mem[12273] = 0;
disk_mem[12274] = 0;
disk_mem[12275] = 0;
disk_mem[12276] = 0;
disk_mem[12277] = 0;
disk_mem[12278] = 0;
disk_mem[12279] = 0;
disk_mem[12280] = 0;
disk_mem[12281] = 0;
disk_mem[12282] = 0;
disk_mem[12283] = 0;
disk_mem[12284] = 0;
disk_mem[12285] = 0;
disk_mem[12286] = 0;
disk_mem[12287] = 0;
disk_mem[12288] = 0;
disk_mem[12289] = 0;
disk_mem[12290] = 0;
disk_mem[12291] = 0;
disk_mem[12292] = 0;
disk_mem[12293] = 0;
disk_mem[12294] = 0;
disk_mem[12295] = 0;
disk_mem[12296] = 0;
disk_mem[12297] = 0;
disk_mem[12298] = 0;
disk_mem[12299] = 0;
disk_mem[12300] = 0;
disk_mem[12301] = 0;
disk_mem[12302] = 0;
disk_mem[12303] = 0;
disk_mem[12304] = 0;
disk_mem[12305] = 0;
disk_mem[12306] = 0;
disk_mem[12307] = 0;
disk_mem[12308] = 0;
disk_mem[12309] = 0;
disk_mem[12310] = 0;
disk_mem[12311] = 0;
disk_mem[12312] = 0;
disk_mem[12313] = 0;
disk_mem[12314] = 0;
disk_mem[12315] = 0;
disk_mem[12316] = 0;
disk_mem[12317] = 0;
disk_mem[12318] = 0;
disk_mem[12319] = 0;
disk_mem[12320] = 0;
disk_mem[12321] = 0;
disk_mem[12322] = 0;
disk_mem[12323] = 0;
disk_mem[12324] = 0;
disk_mem[12325] = 0;
disk_mem[12326] = 0;
disk_mem[12327] = 0;
disk_mem[12328] = 0;
disk_mem[12329] = 0;
disk_mem[12330] = 0;
disk_mem[12331] = 0;
disk_mem[12332] = 0;
disk_mem[12333] = 0;
disk_mem[12334] = 0;
disk_mem[12335] = 0;
disk_mem[12336] = 0;
disk_mem[12337] = 0;
disk_mem[12338] = 0;
disk_mem[12339] = 0;
disk_mem[12340] = 0;
disk_mem[12341] = 0;
disk_mem[12342] = 0;
disk_mem[12343] = 0;
disk_mem[12344] = 0;
disk_mem[12345] = 0;
disk_mem[12346] = 0;
disk_mem[12347] = 0;
disk_mem[12348] = 0;
disk_mem[12349] = 0;
disk_mem[12350] = 0;
disk_mem[12351] = 0;
disk_mem[12352] = 0;
disk_mem[12353] = 0;
disk_mem[12354] = 0;
disk_mem[12355] = 0;
disk_mem[12356] = 0;
disk_mem[12357] = 0;
disk_mem[12358] = 0;
disk_mem[12359] = 0;
disk_mem[12360] = 0;
disk_mem[12361] = 0;
disk_mem[12362] = 0;
disk_mem[12363] = 0;
disk_mem[12364] = 0;
disk_mem[12365] = 0;
disk_mem[12366] = 0;
disk_mem[12367] = 0;
disk_mem[12368] = 0;
disk_mem[12369] = 0;
disk_mem[12370] = 0;
disk_mem[12371] = 0;
disk_mem[12372] = 0;
disk_mem[12373] = 0;
disk_mem[12374] = 0;
disk_mem[12375] = 0;
disk_mem[12376] = 0;
disk_mem[12377] = 0;
disk_mem[12378] = 0;
disk_mem[12379] = 0;
disk_mem[12380] = 0;
disk_mem[12381] = 0;
disk_mem[12382] = 0;
disk_mem[12383] = 0;
disk_mem[12384] = 0;
disk_mem[12385] = 0;
disk_mem[12386] = 0;
disk_mem[12387] = 0;
disk_mem[12388] = 0;
disk_mem[12389] = 0;
disk_mem[12390] = 0;
disk_mem[12391] = 0;
disk_mem[12392] = 0;
disk_mem[12393] = 0;
disk_mem[12394] = 0;
disk_mem[12395] = 0;
disk_mem[12396] = 0;
disk_mem[12397] = 0;
disk_mem[12398] = 0;
disk_mem[12399] = 0;
disk_mem[12400] = 0;
disk_mem[12401] = 0;
disk_mem[12402] = 0;
disk_mem[12403] = 0;
disk_mem[12404] = 0;
disk_mem[12405] = 0;
disk_mem[12406] = 0;
disk_mem[12407] = 0;
disk_mem[12408] = 0;
disk_mem[12409] = 0;
disk_mem[12410] = 0;
disk_mem[12411] = 0;
disk_mem[12412] = 0;
disk_mem[12413] = 0;
disk_mem[12414] = 0;
disk_mem[12415] = 0;
disk_mem[12416] = 0;
disk_mem[12417] = 0;
disk_mem[12418] = 0;
disk_mem[12419] = 0;
disk_mem[12420] = 0;
disk_mem[12421] = 0;
disk_mem[12422] = 0;
disk_mem[12423] = 0;
disk_mem[12424] = 0;
disk_mem[12425] = 0;
disk_mem[12426] = 0;
disk_mem[12427] = 0;
disk_mem[12428] = 0;
disk_mem[12429] = 0;
disk_mem[12430] = 0;
disk_mem[12431] = 0;
disk_mem[12432] = 0;
disk_mem[12433] = 0;
disk_mem[12434] = 0;
disk_mem[12435] = 0;
disk_mem[12436] = 0;
disk_mem[12437] = 0;
disk_mem[12438] = 0;
disk_mem[12439] = 0;
disk_mem[12440] = 0;
disk_mem[12441] = 0;
disk_mem[12442] = 0;
disk_mem[12443] = 0;
disk_mem[12444] = 0;
disk_mem[12445] = 0;
disk_mem[12446] = 0;
disk_mem[12447] = 0;
disk_mem[12448] = 0;
disk_mem[12449] = 0;
disk_mem[12450] = 0;
disk_mem[12451] = 0;
disk_mem[12452] = 0;
disk_mem[12453] = 0;
disk_mem[12454] = 0;
disk_mem[12455] = 0;
disk_mem[12456] = 0;
disk_mem[12457] = 0;
disk_mem[12458] = 0;
disk_mem[12459] = 0;
disk_mem[12460] = 0;
disk_mem[12461] = 0;
disk_mem[12462] = 0;
disk_mem[12463] = 0;
disk_mem[12464] = 0;
disk_mem[12465] = 0;
disk_mem[12466] = 0;
disk_mem[12467] = 0;
disk_mem[12468] = 0;
disk_mem[12469] = 0;
disk_mem[12470] = 0;
disk_mem[12471] = 0;
disk_mem[12472] = 0;
disk_mem[12473] = 0;
disk_mem[12474] = 0;
disk_mem[12475] = 0;
disk_mem[12476] = 0;
disk_mem[12477] = 0;
disk_mem[12478] = 0;
disk_mem[12479] = 0;
disk_mem[12480] = 0;
disk_mem[12481] = 0;
disk_mem[12482] = 0;
disk_mem[12483] = 0;
disk_mem[12484] = 0;
disk_mem[12485] = 0;
disk_mem[12486] = 0;
disk_mem[12487] = 0;
disk_mem[12488] = 0;
disk_mem[12489] = 0;
disk_mem[12490] = 0;
disk_mem[12491] = 0;
disk_mem[12492] = 0;
disk_mem[12493] = 0;
disk_mem[12494] = 0;
disk_mem[12495] = 0;
disk_mem[12496] = 0;
disk_mem[12497] = 0;
disk_mem[12498] = 0;
disk_mem[12499] = 0;
disk_mem[12500] = 0;
disk_mem[12501] = 0;
disk_mem[12502] = 0;
disk_mem[12503] = 0;
disk_mem[12504] = 0;
disk_mem[12505] = 0;
disk_mem[12506] = 0;
disk_mem[12507] = 0;
disk_mem[12508] = 0;
disk_mem[12509] = 0;
disk_mem[12510] = 0;
disk_mem[12511] = 0;
disk_mem[12512] = 0;
disk_mem[12513] = 0;
disk_mem[12514] = 0;
disk_mem[12515] = 0;
disk_mem[12516] = 0;
disk_mem[12517] = 0;
disk_mem[12518] = 0;
disk_mem[12519] = 0;
disk_mem[12520] = 0;
disk_mem[12521] = 0;
disk_mem[12522] = 0;
disk_mem[12523] = 0;
disk_mem[12524] = 0;
disk_mem[12525] = 0;
disk_mem[12526] = 0;
disk_mem[12527] = 0;
disk_mem[12528] = 0;
disk_mem[12529] = 0;
disk_mem[12530] = 0;
disk_mem[12531] = 0;
disk_mem[12532] = 0;
disk_mem[12533] = 0;
disk_mem[12534] = 0;
disk_mem[12535] = 0;
disk_mem[12536] = 0;
disk_mem[12537] = 0;
disk_mem[12538] = 0;
disk_mem[12539] = 0;
disk_mem[12540] = 0;
disk_mem[12541] = 0;
disk_mem[12542] = 0;
disk_mem[12543] = 0;
disk_mem[12544] = 0;
disk_mem[12545] = 0;
disk_mem[12546] = 0;
disk_mem[12547] = 0;
disk_mem[12548] = 0;
disk_mem[12549] = 0;
disk_mem[12550] = 0;
disk_mem[12551] = 0;
disk_mem[12552] = 0;
disk_mem[12553] = 0;
disk_mem[12554] = 0;
disk_mem[12555] = 0;
disk_mem[12556] = 0;
disk_mem[12557] = 0;
disk_mem[12558] = 0;
disk_mem[12559] = 0;
disk_mem[12560] = 0;
disk_mem[12561] = 0;
disk_mem[12562] = 0;
disk_mem[12563] = 0;
disk_mem[12564] = 0;
disk_mem[12565] = 0;
disk_mem[12566] = 0;
disk_mem[12567] = 0;
disk_mem[12568] = 0;
disk_mem[12569] = 0;
disk_mem[12570] = 0;
disk_mem[12571] = 0;
disk_mem[12572] = 0;
disk_mem[12573] = 0;
disk_mem[12574] = 0;
disk_mem[12575] = 0;
disk_mem[12576] = 0;
disk_mem[12577] = 0;
disk_mem[12578] = 0;
disk_mem[12579] = 0;
disk_mem[12580] = 0;
disk_mem[12581] = 0;
disk_mem[12582] = 0;
disk_mem[12583] = 0;
disk_mem[12584] = 0;
disk_mem[12585] = 0;
disk_mem[12586] = 0;
disk_mem[12587] = 0;
disk_mem[12588] = 0;
disk_mem[12589] = 0;
disk_mem[12590] = 0;
disk_mem[12591] = 0;
disk_mem[12592] = 0;
disk_mem[12593] = 0;
disk_mem[12594] = 0;
disk_mem[12595] = 0;
disk_mem[12596] = 0;
disk_mem[12597] = 0;
disk_mem[12598] = 0;
disk_mem[12599] = 0;
disk_mem[12600] = 0;
disk_mem[12601] = 0;
disk_mem[12602] = 0;
disk_mem[12603] = 0;
disk_mem[12604] = 0;
disk_mem[12605] = 0;
disk_mem[12606] = 0;
disk_mem[12607] = 0;
disk_mem[12608] = 0;
disk_mem[12609] = 0;
disk_mem[12610] = 0;
disk_mem[12611] = 0;
disk_mem[12612] = 0;
disk_mem[12613] = 0;
disk_mem[12614] = 0;
disk_mem[12615] = 0;
disk_mem[12616] = 0;
disk_mem[12617] = 0;
disk_mem[12618] = 0;
disk_mem[12619] = 0;
disk_mem[12620] = 0;
disk_mem[12621] = 0;
disk_mem[12622] = 0;
disk_mem[12623] = 0;
disk_mem[12624] = 0;
disk_mem[12625] = 0;
disk_mem[12626] = 0;
disk_mem[12627] = 0;
disk_mem[12628] = 0;
disk_mem[12629] = 0;
disk_mem[12630] = 0;
disk_mem[12631] = 0;
disk_mem[12632] = 0;
disk_mem[12633] = 0;
disk_mem[12634] = 0;
disk_mem[12635] = 0;
disk_mem[12636] = 0;
disk_mem[12637] = 0;
disk_mem[12638] = 0;
disk_mem[12639] = 0;
disk_mem[12640] = 0;
disk_mem[12641] = 0;
disk_mem[12642] = 0;
disk_mem[12643] = 0;
disk_mem[12644] = 0;
disk_mem[12645] = 0;
disk_mem[12646] = 0;
disk_mem[12647] = 0;
disk_mem[12648] = 0;
disk_mem[12649] = 0;
disk_mem[12650] = 0;
disk_mem[12651] = 0;
disk_mem[12652] = 0;
disk_mem[12653] = 0;
disk_mem[12654] = 0;
disk_mem[12655] = 0;
disk_mem[12656] = 0;
disk_mem[12657] = 0;
disk_mem[12658] = 0;
disk_mem[12659] = 0;
disk_mem[12660] = 0;
disk_mem[12661] = 0;
disk_mem[12662] = 0;
disk_mem[12663] = 0;
disk_mem[12664] = 0;
disk_mem[12665] = 0;
disk_mem[12666] = 0;
disk_mem[12667] = 0;
disk_mem[12668] = 0;
disk_mem[12669] = 0;
disk_mem[12670] = 0;
disk_mem[12671] = 0;
disk_mem[12672] = 0;
disk_mem[12673] = 0;
disk_mem[12674] = 0;
disk_mem[12675] = 0;
disk_mem[12676] = 0;
disk_mem[12677] = 0;
disk_mem[12678] = 0;
disk_mem[12679] = 0;
disk_mem[12680] = 0;
disk_mem[12681] = 0;
disk_mem[12682] = 0;
disk_mem[12683] = 0;
disk_mem[12684] = 0;
disk_mem[12685] = 0;
disk_mem[12686] = 0;
disk_mem[12687] = 0;
disk_mem[12688] = 0;
disk_mem[12689] = 0;
disk_mem[12690] = 0;
disk_mem[12691] = 0;
disk_mem[12692] = 0;
disk_mem[12693] = 0;
disk_mem[12694] = 0;
disk_mem[12695] = 0;
disk_mem[12696] = 0;
disk_mem[12697] = 0;
disk_mem[12698] = 0;
disk_mem[12699] = 0;
disk_mem[12700] = 0;
disk_mem[12701] = 0;
disk_mem[12702] = 0;
disk_mem[12703] = 0;
disk_mem[12704] = 0;
disk_mem[12705] = 0;
disk_mem[12706] = 0;
disk_mem[12707] = 0;
disk_mem[12708] = 0;
disk_mem[12709] = 0;
disk_mem[12710] = 0;
disk_mem[12711] = 0;
disk_mem[12712] = 0;
disk_mem[12713] = 0;
disk_mem[12714] = 0;
disk_mem[12715] = 0;
disk_mem[12716] = 0;
disk_mem[12717] = 0;
disk_mem[12718] = 0;
disk_mem[12719] = 0;
disk_mem[12720] = 0;
disk_mem[12721] = 0;
disk_mem[12722] = 0;
disk_mem[12723] = 0;
disk_mem[12724] = 0;
disk_mem[12725] = 0;
disk_mem[12726] = 0;
disk_mem[12727] = 0;
disk_mem[12728] = 0;
disk_mem[12729] = 0;
disk_mem[12730] = 0;
disk_mem[12731] = 0;
disk_mem[12732] = 0;
disk_mem[12733] = 0;
disk_mem[12734] = 0;
disk_mem[12735] = 0;
disk_mem[12736] = 0;
disk_mem[12737] = 0;
disk_mem[12738] = 0;
disk_mem[12739] = 0;
disk_mem[12740] = 0;
disk_mem[12741] = 0;
disk_mem[12742] = 0;
disk_mem[12743] = 0;
disk_mem[12744] = 0;
disk_mem[12745] = 0;
disk_mem[12746] = 0;
disk_mem[12747] = 0;
disk_mem[12748] = 0;
disk_mem[12749] = 0;
disk_mem[12750] = 0;
disk_mem[12751] = 0;
disk_mem[12752] = 0;
disk_mem[12753] = 0;
disk_mem[12754] = 0;
disk_mem[12755] = 0;
disk_mem[12756] = 0;
disk_mem[12757] = 0;
disk_mem[12758] = 0;
disk_mem[12759] = 0;
disk_mem[12760] = 0;
disk_mem[12761] = 0;
disk_mem[12762] = 0;
disk_mem[12763] = 0;
disk_mem[12764] = 0;
disk_mem[12765] = 0;
disk_mem[12766] = 0;
disk_mem[12767] = 0;
disk_mem[12768] = 0;
disk_mem[12769] = 0;
disk_mem[12770] = 0;
disk_mem[12771] = 0;
disk_mem[12772] = 0;
disk_mem[12773] = 0;
disk_mem[12774] = 0;
disk_mem[12775] = 0;
disk_mem[12776] = 0;
disk_mem[12777] = 0;
disk_mem[12778] = 0;
disk_mem[12779] = 0;
disk_mem[12780] = 0;
disk_mem[12781] = 0;
disk_mem[12782] = 0;
disk_mem[12783] = 0;
disk_mem[12784] = 0;
disk_mem[12785] = 0;
disk_mem[12786] = 0;
disk_mem[12787] = 0;
disk_mem[12788] = 0;
disk_mem[12789] = 0;
disk_mem[12790] = 0;
disk_mem[12791] = 0;
disk_mem[12792] = 0;
disk_mem[12793] = 0;
disk_mem[12794] = 0;
disk_mem[12795] = 0;
disk_mem[12796] = 0;
disk_mem[12797] = 0;
disk_mem[12798] = 0;
disk_mem[12799] = 0;
disk_mem[12800] = 0;
disk_mem[12801] = 0;
disk_mem[12802] = 0;
disk_mem[12803] = 0;
disk_mem[12804] = 0;
disk_mem[12805] = 0;
disk_mem[12806] = 0;
disk_mem[12807] = 0;
disk_mem[12808] = 0;
disk_mem[12809] = 0;
disk_mem[12810] = 0;
disk_mem[12811] = 0;
disk_mem[12812] = 0;
disk_mem[12813] = 0;
disk_mem[12814] = 0;
disk_mem[12815] = 0;
disk_mem[12816] = 0;
disk_mem[12817] = 0;
disk_mem[12818] = 0;
disk_mem[12819] = 0;
disk_mem[12820] = 0;
disk_mem[12821] = 0;
disk_mem[12822] = 0;
disk_mem[12823] = 0;
disk_mem[12824] = 0;
disk_mem[12825] = 0;
disk_mem[12826] = 0;
disk_mem[12827] = 0;
disk_mem[12828] = 0;
disk_mem[12829] = 0;
disk_mem[12830] = 0;
disk_mem[12831] = 0;
disk_mem[12832] = 0;
disk_mem[12833] = 0;
disk_mem[12834] = 0;
disk_mem[12835] = 0;
disk_mem[12836] = 0;
disk_mem[12837] = 0;
disk_mem[12838] = 0;
disk_mem[12839] = 0;
disk_mem[12840] = 0;
disk_mem[12841] = 0;
disk_mem[12842] = 0;
disk_mem[12843] = 0;
disk_mem[12844] = 0;
disk_mem[12845] = 0;
disk_mem[12846] = 0;
disk_mem[12847] = 0;
disk_mem[12848] = 0;
disk_mem[12849] = 0;
disk_mem[12850] = 0;
disk_mem[12851] = 0;
disk_mem[12852] = 0;
disk_mem[12853] = 0;
disk_mem[12854] = 0;
disk_mem[12855] = 0;
disk_mem[12856] = 0;
disk_mem[12857] = 0;
disk_mem[12858] = 0;
disk_mem[12859] = 0;
disk_mem[12860] = 0;
disk_mem[12861] = 0;
disk_mem[12862] = 0;
disk_mem[12863] = 0;
disk_mem[12864] = 0;
disk_mem[12865] = 0;
disk_mem[12866] = 0;
disk_mem[12867] = 0;
disk_mem[12868] = 0;
disk_mem[12869] = 0;
disk_mem[12870] = 0;
disk_mem[12871] = 0;
disk_mem[12872] = 0;
disk_mem[12873] = 0;
disk_mem[12874] = 0;
disk_mem[12875] = 0;
disk_mem[12876] = 0;
disk_mem[12877] = 0;
disk_mem[12878] = 0;
disk_mem[12879] = 0;
disk_mem[12880] = 0;
disk_mem[12881] = 0;
disk_mem[12882] = 0;
disk_mem[12883] = 0;
disk_mem[12884] = 0;
disk_mem[12885] = 0;
disk_mem[12886] = 0;
disk_mem[12887] = 0;
disk_mem[12888] = 0;
disk_mem[12889] = 0;
disk_mem[12890] = 0;
disk_mem[12891] = 0;
disk_mem[12892] = 0;
disk_mem[12893] = 0;
disk_mem[12894] = 0;
disk_mem[12895] = 0;
disk_mem[12896] = 0;
disk_mem[12897] = 0;
disk_mem[12898] = 0;
disk_mem[12899] = 0;
disk_mem[12900] = 0;
disk_mem[12901] = 0;
disk_mem[12902] = 0;
disk_mem[12903] = 0;
disk_mem[12904] = 0;
disk_mem[12905] = 0;
disk_mem[12906] = 0;
disk_mem[12907] = 0;
disk_mem[12908] = 0;
disk_mem[12909] = 0;
disk_mem[12910] = 0;
disk_mem[12911] = 0;
disk_mem[12912] = 0;
disk_mem[12913] = 0;
disk_mem[12914] = 0;
disk_mem[12915] = 0;
disk_mem[12916] = 0;
disk_mem[12917] = 0;
disk_mem[12918] = 0;
disk_mem[12919] = 0;
disk_mem[12920] = 0;
disk_mem[12921] = 0;
disk_mem[12922] = 0;
disk_mem[12923] = 0;
disk_mem[12924] = 0;
disk_mem[12925] = 0;
disk_mem[12926] = 0;
disk_mem[12927] = 0;
disk_mem[12928] = 0;
disk_mem[12929] = 0;
disk_mem[12930] = 0;
disk_mem[12931] = 0;
disk_mem[12932] = 0;
disk_mem[12933] = 0;
disk_mem[12934] = 0;
disk_mem[12935] = 0;
disk_mem[12936] = 0;
disk_mem[12937] = 0;
disk_mem[12938] = 0;
disk_mem[12939] = 0;
disk_mem[12940] = 0;
disk_mem[12941] = 0;
disk_mem[12942] = 0;
disk_mem[12943] = 0;
disk_mem[12944] = 0;
disk_mem[12945] = 0;
disk_mem[12946] = 0;
disk_mem[12947] = 0;
disk_mem[12948] = 0;
disk_mem[12949] = 0;
disk_mem[12950] = 0;
disk_mem[12951] = 0;
disk_mem[12952] = 0;
disk_mem[12953] = 0;
disk_mem[12954] = 0;
disk_mem[12955] = 0;
disk_mem[12956] = 0;
disk_mem[12957] = 0;
disk_mem[12958] = 0;
disk_mem[12959] = 0;
disk_mem[12960] = 0;
disk_mem[12961] = 0;
disk_mem[12962] = 0;
disk_mem[12963] = 0;
disk_mem[12964] = 0;
disk_mem[12965] = 0;
disk_mem[12966] = 0;
disk_mem[12967] = 0;
disk_mem[12968] = 0;
disk_mem[12969] = 0;
disk_mem[12970] = 0;
disk_mem[12971] = 0;
disk_mem[12972] = 0;
disk_mem[12973] = 0;
disk_mem[12974] = 0;
disk_mem[12975] = 0;
disk_mem[12976] = 0;
disk_mem[12977] = 0;
disk_mem[12978] = 0;
disk_mem[12979] = 0;
disk_mem[12980] = 0;
disk_mem[12981] = 0;
disk_mem[12982] = 0;
disk_mem[12983] = 0;
disk_mem[12984] = 0;
disk_mem[12985] = 0;
disk_mem[12986] = 0;
disk_mem[12987] = 0;
disk_mem[12988] = 0;
disk_mem[12989] = 0;
disk_mem[12990] = 0;
disk_mem[12991] = 0;
disk_mem[12992] = 0;
disk_mem[12993] = 0;
disk_mem[12994] = 0;
disk_mem[12995] = 0;
disk_mem[12996] = 0;
disk_mem[12997] = 0;
disk_mem[12998] = 0;
disk_mem[12999] = 0;
disk_mem[13000] = 0;
disk_mem[13001] = 0;
disk_mem[13002] = 0;
disk_mem[13003] = 0;
disk_mem[13004] = 0;
disk_mem[13005] = 0;
disk_mem[13006] = 0;
disk_mem[13007] = 0;
disk_mem[13008] = 0;
disk_mem[13009] = 0;
disk_mem[13010] = 0;
disk_mem[13011] = 0;
disk_mem[13012] = 0;
disk_mem[13013] = 0;
disk_mem[13014] = 0;
disk_mem[13015] = 0;
disk_mem[13016] = 0;
disk_mem[13017] = 0;
disk_mem[13018] = 0;
disk_mem[13019] = 0;
disk_mem[13020] = 0;
disk_mem[13021] = 0;
disk_mem[13022] = 0;
disk_mem[13023] = 0;
disk_mem[13024] = 0;
disk_mem[13025] = 0;
disk_mem[13026] = 0;
disk_mem[13027] = 0;
disk_mem[13028] = 0;
disk_mem[13029] = 0;
disk_mem[13030] = 0;
disk_mem[13031] = 0;
disk_mem[13032] = 0;
disk_mem[13033] = 0;
disk_mem[13034] = 0;
disk_mem[13035] = 0;
disk_mem[13036] = 0;
disk_mem[13037] = 0;
disk_mem[13038] = 0;
disk_mem[13039] = 0;
disk_mem[13040] = 0;
disk_mem[13041] = 0;
disk_mem[13042] = 0;
disk_mem[13043] = 0;
disk_mem[13044] = 0;
disk_mem[13045] = 0;
disk_mem[13046] = 0;
disk_mem[13047] = 0;
disk_mem[13048] = 0;
disk_mem[13049] = 0;
disk_mem[13050] = 0;
disk_mem[13051] = 0;
disk_mem[13052] = 0;
disk_mem[13053] = 0;
disk_mem[13054] = 0;
disk_mem[13055] = 0;
disk_mem[13056] = 0;
disk_mem[13057] = 0;
disk_mem[13058] = 0;
disk_mem[13059] = 0;
disk_mem[13060] = 0;
disk_mem[13061] = 0;
disk_mem[13062] = 0;
disk_mem[13063] = 0;
disk_mem[13064] = 0;
disk_mem[13065] = 0;
disk_mem[13066] = 0;
disk_mem[13067] = 0;
disk_mem[13068] = 0;
disk_mem[13069] = 0;
disk_mem[13070] = 0;
disk_mem[13071] = 0;
disk_mem[13072] = 0;
disk_mem[13073] = 0;
disk_mem[13074] = 0;
disk_mem[13075] = 0;
disk_mem[13076] = 0;
disk_mem[13077] = 0;
disk_mem[13078] = 0;
disk_mem[13079] = 0;
disk_mem[13080] = 0;
disk_mem[13081] = 0;
disk_mem[13082] = 0;
disk_mem[13083] = 0;
disk_mem[13084] = 0;
disk_mem[13085] = 0;
disk_mem[13086] = 0;
disk_mem[13087] = 0;
disk_mem[13088] = 0;
disk_mem[13089] = 0;
disk_mem[13090] = 0;
disk_mem[13091] = 0;
disk_mem[13092] = 0;
disk_mem[13093] = 0;
disk_mem[13094] = 0;
disk_mem[13095] = 0;
disk_mem[13096] = 0;
disk_mem[13097] = 0;
disk_mem[13098] = 0;
disk_mem[13099] = 0;
disk_mem[13100] = 0;
disk_mem[13101] = 0;
disk_mem[13102] = 0;
disk_mem[13103] = 0;
disk_mem[13104] = 0;
disk_mem[13105] = 0;
disk_mem[13106] = 0;
disk_mem[13107] = 0;
disk_mem[13108] = 0;
disk_mem[13109] = 0;
disk_mem[13110] = 0;
disk_mem[13111] = 0;
disk_mem[13112] = 0;
disk_mem[13113] = 0;
disk_mem[13114] = 0;
disk_mem[13115] = 0;
disk_mem[13116] = 0;
disk_mem[13117] = 0;
disk_mem[13118] = 0;
disk_mem[13119] = 0;
disk_mem[13120] = 0;
disk_mem[13121] = 0;
disk_mem[13122] = 0;
disk_mem[13123] = 0;
disk_mem[13124] = 0;
disk_mem[13125] = 0;
disk_mem[13126] = 0;
disk_mem[13127] = 0;
disk_mem[13128] = 0;
disk_mem[13129] = 0;
disk_mem[13130] = 0;
disk_mem[13131] = 0;
disk_mem[13132] = 0;
disk_mem[13133] = 0;
disk_mem[13134] = 0;
disk_mem[13135] = 0;
disk_mem[13136] = 0;
disk_mem[13137] = 0;
disk_mem[13138] = 0;
disk_mem[13139] = 0;
disk_mem[13140] = 0;
disk_mem[13141] = 0;
disk_mem[13142] = 0;
disk_mem[13143] = 0;
disk_mem[13144] = 0;
disk_mem[13145] = 0;
disk_mem[13146] = 0;
disk_mem[13147] = 0;
disk_mem[13148] = 0;
disk_mem[13149] = 0;
disk_mem[13150] = 0;
disk_mem[13151] = 0;
disk_mem[13152] = 0;
disk_mem[13153] = 0;
disk_mem[13154] = 0;
disk_mem[13155] = 0;
disk_mem[13156] = 0;
disk_mem[13157] = 0;
disk_mem[13158] = 0;
disk_mem[13159] = 0;
disk_mem[13160] = 0;
disk_mem[13161] = 0;
disk_mem[13162] = 0;
disk_mem[13163] = 0;
disk_mem[13164] = 0;
disk_mem[13165] = 0;
disk_mem[13166] = 0;
disk_mem[13167] = 0;
disk_mem[13168] = 0;
disk_mem[13169] = 0;
disk_mem[13170] = 0;
disk_mem[13171] = 0;
disk_mem[13172] = 0;
disk_mem[13173] = 0;
disk_mem[13174] = 0;
disk_mem[13175] = 0;
disk_mem[13176] = 0;
disk_mem[13177] = 0;
disk_mem[13178] = 0;
disk_mem[13179] = 0;
disk_mem[13180] = 0;
disk_mem[13181] = 0;
disk_mem[13182] = 0;
disk_mem[13183] = 0;
disk_mem[13184] = 0;
disk_mem[13185] = 0;
disk_mem[13186] = 0;
disk_mem[13187] = 0;
disk_mem[13188] = 0;
disk_mem[13189] = 0;
disk_mem[13190] = 0;
disk_mem[13191] = 0;
disk_mem[13192] = 0;
disk_mem[13193] = 0;
disk_mem[13194] = 0;
disk_mem[13195] = 0;
disk_mem[13196] = 0;
disk_mem[13197] = 0;
disk_mem[13198] = 0;
disk_mem[13199] = 0;
disk_mem[13200] = 0;
disk_mem[13201] = 0;
disk_mem[13202] = 0;
disk_mem[13203] = 0;
disk_mem[13204] = 0;
disk_mem[13205] = 0;
disk_mem[13206] = 0;
disk_mem[13207] = 0;
disk_mem[13208] = 0;
disk_mem[13209] = 0;
disk_mem[13210] = 0;
disk_mem[13211] = 0;
disk_mem[13212] = 0;
disk_mem[13213] = 0;
disk_mem[13214] = 0;
disk_mem[13215] = 0;
disk_mem[13216] = 0;
disk_mem[13217] = 0;
disk_mem[13218] = 0;
disk_mem[13219] = 0;
disk_mem[13220] = 0;
disk_mem[13221] = 0;
disk_mem[13222] = 0;
disk_mem[13223] = 0;
disk_mem[13224] = 0;
disk_mem[13225] = 0;
disk_mem[13226] = 0;
disk_mem[13227] = 0;
disk_mem[13228] = 0;
disk_mem[13229] = 0;
disk_mem[13230] = 0;
disk_mem[13231] = 0;
disk_mem[13232] = 0;
disk_mem[13233] = 0;
disk_mem[13234] = 0;
disk_mem[13235] = 0;
disk_mem[13236] = 0;
disk_mem[13237] = 0;
disk_mem[13238] = 0;
disk_mem[13239] = 0;
disk_mem[13240] = 0;
disk_mem[13241] = 0;
disk_mem[13242] = 0;
disk_mem[13243] = 0;
disk_mem[13244] = 0;
disk_mem[13245] = 0;
disk_mem[13246] = 0;
disk_mem[13247] = 0;
disk_mem[13248] = 0;
disk_mem[13249] = 0;
disk_mem[13250] = 0;
disk_mem[13251] = 0;
disk_mem[13252] = 0;
disk_mem[13253] = 0;
disk_mem[13254] = 0;
disk_mem[13255] = 0;
disk_mem[13256] = 0;
disk_mem[13257] = 0;
disk_mem[13258] = 0;
disk_mem[13259] = 0;
disk_mem[13260] = 0;
disk_mem[13261] = 0;
disk_mem[13262] = 0;
disk_mem[13263] = 0;
disk_mem[13264] = 0;
disk_mem[13265] = 0;
disk_mem[13266] = 0;
disk_mem[13267] = 0;
disk_mem[13268] = 0;
disk_mem[13269] = 0;
disk_mem[13270] = 0;
disk_mem[13271] = 0;
disk_mem[13272] = 0;
disk_mem[13273] = 0;
disk_mem[13274] = 0;
disk_mem[13275] = 0;
disk_mem[13276] = 0;
disk_mem[13277] = 0;
disk_mem[13278] = 0;
disk_mem[13279] = 0;
disk_mem[13280] = 0;
disk_mem[13281] = 0;
disk_mem[13282] = 0;
disk_mem[13283] = 0;
disk_mem[13284] = 0;
disk_mem[13285] = 0;
disk_mem[13286] = 0;
disk_mem[13287] = 0;
disk_mem[13288] = 0;
disk_mem[13289] = 0;
disk_mem[13290] = 0;
disk_mem[13291] = 0;
disk_mem[13292] = 0;
disk_mem[13293] = 0;
disk_mem[13294] = 0;
disk_mem[13295] = 0;
disk_mem[13296] = 0;
disk_mem[13297] = 0;
disk_mem[13298] = 0;
disk_mem[13299] = 0;
disk_mem[13300] = 0;
disk_mem[13301] = 0;
disk_mem[13302] = 0;
disk_mem[13303] = 0;
disk_mem[13304] = 0;
disk_mem[13305] = 0;
disk_mem[13306] = 0;
disk_mem[13307] = 0;
disk_mem[13308] = 0;
disk_mem[13309] = 0;
disk_mem[13310] = 0;
disk_mem[13311] = 0;
disk_mem[13312] = 0;
disk_mem[13313] = 0;
disk_mem[13314] = 0;
disk_mem[13315] = 0;
disk_mem[13316] = 0;
disk_mem[13317] = 0;
disk_mem[13318] = 0;
disk_mem[13319] = 0;
disk_mem[13320] = 0;
disk_mem[13321] = 0;
disk_mem[13322] = 0;
disk_mem[13323] = 0;
disk_mem[13324] = 0;
disk_mem[13325] = 0;
disk_mem[13326] = 0;
disk_mem[13327] = 0;
disk_mem[13328] = 0;
disk_mem[13329] = 0;
disk_mem[13330] = 0;
disk_mem[13331] = 0;
disk_mem[13332] = 0;
disk_mem[13333] = 0;
disk_mem[13334] = 0;
disk_mem[13335] = 0;
disk_mem[13336] = 0;
disk_mem[13337] = 0;
disk_mem[13338] = 0;
disk_mem[13339] = 0;
disk_mem[13340] = 0;
disk_mem[13341] = 0;
disk_mem[13342] = 0;
disk_mem[13343] = 0;
disk_mem[13344] = 0;
disk_mem[13345] = 0;
disk_mem[13346] = 0;
disk_mem[13347] = 0;
disk_mem[13348] = 0;
disk_mem[13349] = 0;
disk_mem[13350] = 0;
disk_mem[13351] = 0;
disk_mem[13352] = 0;
disk_mem[13353] = 0;
disk_mem[13354] = 0;
disk_mem[13355] = 0;
disk_mem[13356] = 0;
disk_mem[13357] = 0;
disk_mem[13358] = 0;
disk_mem[13359] = 0;
disk_mem[13360] = 0;
disk_mem[13361] = 0;
disk_mem[13362] = 0;
disk_mem[13363] = 0;
disk_mem[13364] = 0;
disk_mem[13365] = 0;
disk_mem[13366] = 0;
disk_mem[13367] = 0;
disk_mem[13368] = 0;
disk_mem[13369] = 0;
disk_mem[13370] = 0;
disk_mem[13371] = 0;
disk_mem[13372] = 0;
disk_mem[13373] = 0;
disk_mem[13374] = 0;
disk_mem[13375] = 0;
disk_mem[13376] = 0;
disk_mem[13377] = 0;
disk_mem[13378] = 0;
disk_mem[13379] = 0;
disk_mem[13380] = 0;
disk_mem[13381] = 0;
disk_mem[13382] = 0;
disk_mem[13383] = 0;
disk_mem[13384] = 0;
disk_mem[13385] = 0;
disk_mem[13386] = 0;
disk_mem[13387] = 0;
disk_mem[13388] = 0;
disk_mem[13389] = 0;
disk_mem[13390] = 0;
disk_mem[13391] = 0;
disk_mem[13392] = 0;
disk_mem[13393] = 0;
disk_mem[13394] = 0;
disk_mem[13395] = 0;
disk_mem[13396] = 0;
disk_mem[13397] = 0;
disk_mem[13398] = 0;
disk_mem[13399] = 0;
disk_mem[13400] = 0;
disk_mem[13401] = 0;
disk_mem[13402] = 0;
disk_mem[13403] = 0;
disk_mem[13404] = 0;
disk_mem[13405] = 0;
disk_mem[13406] = 0;
disk_mem[13407] = 0;
disk_mem[13408] = 0;
disk_mem[13409] = 0;
disk_mem[13410] = 0;
disk_mem[13411] = 0;
disk_mem[13412] = 0;
disk_mem[13413] = 0;
disk_mem[13414] = 0;
disk_mem[13415] = 0;
disk_mem[13416] = 0;
disk_mem[13417] = 0;
disk_mem[13418] = 0;
disk_mem[13419] = 0;
disk_mem[13420] = 0;
disk_mem[13421] = 0;
disk_mem[13422] = 0;
disk_mem[13423] = 0;
disk_mem[13424] = 0;
disk_mem[13425] = 0;
disk_mem[13426] = 0;
disk_mem[13427] = 0;
disk_mem[13428] = 0;
disk_mem[13429] = 0;
disk_mem[13430] = 0;
disk_mem[13431] = 0;
disk_mem[13432] = 0;
disk_mem[13433] = 0;
disk_mem[13434] = 0;
disk_mem[13435] = 0;
disk_mem[13436] = 0;
disk_mem[13437] = 0;
disk_mem[13438] = 0;
disk_mem[13439] = 0;
disk_mem[13440] = 0;
disk_mem[13441] = 0;
disk_mem[13442] = 0;
disk_mem[13443] = 0;
disk_mem[13444] = 0;
disk_mem[13445] = 0;
disk_mem[13446] = 0;
disk_mem[13447] = 0;
disk_mem[13448] = 0;
disk_mem[13449] = 0;
disk_mem[13450] = 0;
disk_mem[13451] = 0;
disk_mem[13452] = 0;
disk_mem[13453] = 0;
disk_mem[13454] = 0;
disk_mem[13455] = 0;
disk_mem[13456] = 0;
disk_mem[13457] = 0;
disk_mem[13458] = 0;
disk_mem[13459] = 0;
disk_mem[13460] = 0;
disk_mem[13461] = 0;
disk_mem[13462] = 0;
disk_mem[13463] = 0;
disk_mem[13464] = 0;
disk_mem[13465] = 0;
disk_mem[13466] = 0;
disk_mem[13467] = 0;
disk_mem[13468] = 0;
disk_mem[13469] = 0;
disk_mem[13470] = 0;
disk_mem[13471] = 0;
disk_mem[13472] = 0;
disk_mem[13473] = 0;
disk_mem[13474] = 0;
disk_mem[13475] = 0;
disk_mem[13476] = 0;
disk_mem[13477] = 0;
disk_mem[13478] = 0;
disk_mem[13479] = 0;
disk_mem[13480] = 0;
disk_mem[13481] = 0;
disk_mem[13482] = 0;
disk_mem[13483] = 0;
disk_mem[13484] = 0;
disk_mem[13485] = 0;
disk_mem[13486] = 0;
disk_mem[13487] = 0;
disk_mem[13488] = 0;
disk_mem[13489] = 0;
disk_mem[13490] = 0;
disk_mem[13491] = 0;
disk_mem[13492] = 0;
disk_mem[13493] = 0;
disk_mem[13494] = 0;
disk_mem[13495] = 0;
disk_mem[13496] = 0;
disk_mem[13497] = 0;
disk_mem[13498] = 0;
disk_mem[13499] = 0;
disk_mem[13500] = 0;
disk_mem[13501] = 0;
disk_mem[13502] = 0;
disk_mem[13503] = 0;
disk_mem[13504] = 0;
disk_mem[13505] = 0;
disk_mem[13506] = 0;
disk_mem[13507] = 0;
disk_mem[13508] = 0;
disk_mem[13509] = 0;
disk_mem[13510] = 0;
disk_mem[13511] = 0;
disk_mem[13512] = 0;
disk_mem[13513] = 0;
disk_mem[13514] = 0;
disk_mem[13515] = 0;
disk_mem[13516] = 0;
disk_mem[13517] = 0;
disk_mem[13518] = 0;
disk_mem[13519] = 0;
disk_mem[13520] = 0;
disk_mem[13521] = 0;
disk_mem[13522] = 0;
disk_mem[13523] = 0;
disk_mem[13524] = 0;
disk_mem[13525] = 0;
disk_mem[13526] = 0;
disk_mem[13527] = 0;
disk_mem[13528] = 0;
disk_mem[13529] = 0;
disk_mem[13530] = 0;
disk_mem[13531] = 0;
disk_mem[13532] = 0;
disk_mem[13533] = 0;
disk_mem[13534] = 0;
disk_mem[13535] = 0;
disk_mem[13536] = 0;
disk_mem[13537] = 0;
disk_mem[13538] = 0;
disk_mem[13539] = 0;
disk_mem[13540] = 0;
disk_mem[13541] = 0;
disk_mem[13542] = 0;
disk_mem[13543] = 0;
disk_mem[13544] = 0;
disk_mem[13545] = 0;
disk_mem[13546] = 0;
disk_mem[13547] = 0;
disk_mem[13548] = 0;
disk_mem[13549] = 0;
disk_mem[13550] = 0;
disk_mem[13551] = 0;
disk_mem[13552] = 0;
disk_mem[13553] = 0;
disk_mem[13554] = 0;
disk_mem[13555] = 0;
disk_mem[13556] = 0;
disk_mem[13557] = 0;
disk_mem[13558] = 0;
disk_mem[13559] = 0;
disk_mem[13560] = 0;
disk_mem[13561] = 0;
disk_mem[13562] = 0;
disk_mem[13563] = 0;
disk_mem[13564] = 0;
disk_mem[13565] = 0;
disk_mem[13566] = 0;
disk_mem[13567] = 0;
disk_mem[13568] = 0;
disk_mem[13569] = 0;
disk_mem[13570] = 0;
disk_mem[13571] = 0;
disk_mem[13572] = 0;
disk_mem[13573] = 0;
disk_mem[13574] = 0;
disk_mem[13575] = 0;
disk_mem[13576] = 0;
disk_mem[13577] = 0;
disk_mem[13578] = 0;
disk_mem[13579] = 0;
disk_mem[13580] = 0;
disk_mem[13581] = 0;
disk_mem[13582] = 0;
disk_mem[13583] = 0;
disk_mem[13584] = 0;
disk_mem[13585] = 0;
disk_mem[13586] = 0;
disk_mem[13587] = 0;
disk_mem[13588] = 0;
disk_mem[13589] = 0;
disk_mem[13590] = 0;
disk_mem[13591] = 0;
disk_mem[13592] = 0;
disk_mem[13593] = 0;
disk_mem[13594] = 0;
disk_mem[13595] = 0;
disk_mem[13596] = 0;
disk_mem[13597] = 0;
disk_mem[13598] = 0;
disk_mem[13599] = 0;
disk_mem[13600] = 0;
disk_mem[13601] = 0;
disk_mem[13602] = 0;
disk_mem[13603] = 0;
disk_mem[13604] = 0;
disk_mem[13605] = 0;
disk_mem[13606] = 0;
disk_mem[13607] = 0;
disk_mem[13608] = 0;
disk_mem[13609] = 0;
disk_mem[13610] = 0;
disk_mem[13611] = 0;
disk_mem[13612] = 0;
disk_mem[13613] = 0;
disk_mem[13614] = 0;
disk_mem[13615] = 0;
disk_mem[13616] = 0;
disk_mem[13617] = 0;
disk_mem[13618] = 0;
disk_mem[13619] = 0;
disk_mem[13620] = 0;
disk_mem[13621] = 0;
disk_mem[13622] = 0;
disk_mem[13623] = 0;
disk_mem[13624] = 0;
disk_mem[13625] = 0;
disk_mem[13626] = 0;
disk_mem[13627] = 0;
disk_mem[13628] = 0;
disk_mem[13629] = 0;
disk_mem[13630] = 0;
disk_mem[13631] = 0;
disk_mem[13632] = 0;
disk_mem[13633] = 0;
disk_mem[13634] = 0;
disk_mem[13635] = 0;
disk_mem[13636] = 0;
disk_mem[13637] = 0;
disk_mem[13638] = 0;
disk_mem[13639] = 0;
disk_mem[13640] = 0;
disk_mem[13641] = 0;
disk_mem[13642] = 0;
disk_mem[13643] = 0;
disk_mem[13644] = 0;
disk_mem[13645] = 0;
disk_mem[13646] = 0;
disk_mem[13647] = 0;
disk_mem[13648] = 0;
disk_mem[13649] = 0;
disk_mem[13650] = 0;
disk_mem[13651] = 0;
disk_mem[13652] = 0;
disk_mem[13653] = 0;
disk_mem[13654] = 0;
disk_mem[13655] = 0;
disk_mem[13656] = 0;
disk_mem[13657] = 0;
disk_mem[13658] = 0;
disk_mem[13659] = 0;
disk_mem[13660] = 0;
disk_mem[13661] = 0;
disk_mem[13662] = 0;
disk_mem[13663] = 0;
disk_mem[13664] = 0;
disk_mem[13665] = 0;
disk_mem[13666] = 0;
disk_mem[13667] = 0;
disk_mem[13668] = 0;
disk_mem[13669] = 0;
disk_mem[13670] = 0;
disk_mem[13671] = 0;
disk_mem[13672] = 0;
disk_mem[13673] = 0;
disk_mem[13674] = 0;
disk_mem[13675] = 0;
disk_mem[13676] = 0;
disk_mem[13677] = 0;
disk_mem[13678] = 0;
disk_mem[13679] = 0;
disk_mem[13680] = 0;
disk_mem[13681] = 0;
disk_mem[13682] = 0;
disk_mem[13683] = 0;
disk_mem[13684] = 0;
disk_mem[13685] = 0;
disk_mem[13686] = 0;
disk_mem[13687] = 0;
disk_mem[13688] = 0;
disk_mem[13689] = 0;
disk_mem[13690] = 0;
disk_mem[13691] = 0;
disk_mem[13692] = 0;
disk_mem[13693] = 0;
disk_mem[13694] = 0;
disk_mem[13695] = 0;
disk_mem[13696] = 0;
disk_mem[13697] = 0;
disk_mem[13698] = 0;
disk_mem[13699] = 0;
disk_mem[13700] = 0;
disk_mem[13701] = 0;
disk_mem[13702] = 0;
disk_mem[13703] = 0;
disk_mem[13704] = 0;
disk_mem[13705] = 0;
disk_mem[13706] = 0;
disk_mem[13707] = 0;
disk_mem[13708] = 0;
disk_mem[13709] = 0;
disk_mem[13710] = 0;
disk_mem[13711] = 0;
disk_mem[13712] = 0;
disk_mem[13713] = 0;
disk_mem[13714] = 0;
disk_mem[13715] = 0;
disk_mem[13716] = 0;
disk_mem[13717] = 0;
disk_mem[13718] = 0;
disk_mem[13719] = 0;
disk_mem[13720] = 0;
disk_mem[13721] = 0;
disk_mem[13722] = 0;
disk_mem[13723] = 0;
disk_mem[13724] = 0;
disk_mem[13725] = 0;
disk_mem[13726] = 0;
disk_mem[13727] = 0;
disk_mem[13728] = 0;
disk_mem[13729] = 0;
disk_mem[13730] = 0;
disk_mem[13731] = 0;
disk_mem[13732] = 0;
disk_mem[13733] = 0;
disk_mem[13734] = 0;
disk_mem[13735] = 0;
disk_mem[13736] = 0;
disk_mem[13737] = 0;
disk_mem[13738] = 0;
disk_mem[13739] = 0;
disk_mem[13740] = 0;
disk_mem[13741] = 0;
disk_mem[13742] = 0;
disk_mem[13743] = 0;
disk_mem[13744] = 0;
disk_mem[13745] = 0;
disk_mem[13746] = 0;
disk_mem[13747] = 0;
disk_mem[13748] = 0;
disk_mem[13749] = 0;
disk_mem[13750] = 0;
disk_mem[13751] = 0;
disk_mem[13752] = 0;
disk_mem[13753] = 0;
disk_mem[13754] = 0;
disk_mem[13755] = 0;
disk_mem[13756] = 0;
disk_mem[13757] = 0;
disk_mem[13758] = 0;
disk_mem[13759] = 0;
disk_mem[13760] = 0;
disk_mem[13761] = 0;
disk_mem[13762] = 0;
disk_mem[13763] = 0;
disk_mem[13764] = 0;
disk_mem[13765] = 0;
disk_mem[13766] = 0;
disk_mem[13767] = 0;
disk_mem[13768] = 0;
disk_mem[13769] = 0;
disk_mem[13770] = 0;
disk_mem[13771] = 0;
disk_mem[13772] = 0;
disk_mem[13773] = 0;
disk_mem[13774] = 0;
disk_mem[13775] = 0;
disk_mem[13776] = 0;
disk_mem[13777] = 0;
disk_mem[13778] = 0;
disk_mem[13779] = 0;
disk_mem[13780] = 0;
disk_mem[13781] = 0;
disk_mem[13782] = 0;
disk_mem[13783] = 0;
disk_mem[13784] = 0;
disk_mem[13785] = 0;
disk_mem[13786] = 0;
disk_mem[13787] = 0;
disk_mem[13788] = 0;
disk_mem[13789] = 0;
disk_mem[13790] = 0;
disk_mem[13791] = 0;
disk_mem[13792] = 0;
disk_mem[13793] = 0;
disk_mem[13794] = 0;
disk_mem[13795] = 0;
disk_mem[13796] = 0;
disk_mem[13797] = 0;
disk_mem[13798] = 0;
disk_mem[13799] = 0;
disk_mem[13800] = 0;
disk_mem[13801] = 0;
disk_mem[13802] = 0;
disk_mem[13803] = 0;
disk_mem[13804] = 0;
disk_mem[13805] = 0;
disk_mem[13806] = 0;
disk_mem[13807] = 0;
disk_mem[13808] = 0;
disk_mem[13809] = 0;
disk_mem[13810] = 0;
disk_mem[13811] = 0;
disk_mem[13812] = 0;
disk_mem[13813] = 0;
disk_mem[13814] = 0;
disk_mem[13815] = 0;
disk_mem[13816] = 0;
disk_mem[13817] = 0;
disk_mem[13818] = 0;
disk_mem[13819] = 0;
disk_mem[13820] = 0;
disk_mem[13821] = 0;
disk_mem[13822] = 0;
disk_mem[13823] = 0;
disk_mem[13824] = 0;
disk_mem[13825] = 0;
disk_mem[13826] = 0;
disk_mem[13827] = 0;
disk_mem[13828] = 0;
disk_mem[13829] = 0;
disk_mem[13830] = 0;
disk_mem[13831] = 0;
disk_mem[13832] = 0;
disk_mem[13833] = 0;
disk_mem[13834] = 0;
disk_mem[13835] = 0;
disk_mem[13836] = 0;
disk_mem[13837] = 0;
disk_mem[13838] = 0;
disk_mem[13839] = 0;
disk_mem[13840] = 0;
disk_mem[13841] = 0;
disk_mem[13842] = 0;
disk_mem[13843] = 0;
disk_mem[13844] = 0;
disk_mem[13845] = 0;
disk_mem[13846] = 0;
disk_mem[13847] = 0;
disk_mem[13848] = 0;
disk_mem[13849] = 0;
disk_mem[13850] = 0;
disk_mem[13851] = 0;
disk_mem[13852] = 0;
disk_mem[13853] = 0;
disk_mem[13854] = 0;
disk_mem[13855] = 0;
disk_mem[13856] = 0;
disk_mem[13857] = 0;
disk_mem[13858] = 0;
disk_mem[13859] = 0;
disk_mem[13860] = 0;
disk_mem[13861] = 0;
disk_mem[13862] = 0;
disk_mem[13863] = 0;
disk_mem[13864] = 0;
disk_mem[13865] = 0;
disk_mem[13866] = 0;
disk_mem[13867] = 0;
disk_mem[13868] = 0;
disk_mem[13869] = 0;
disk_mem[13870] = 0;
disk_mem[13871] = 0;
disk_mem[13872] = 0;
disk_mem[13873] = 0;
disk_mem[13874] = 0;
disk_mem[13875] = 0;
disk_mem[13876] = 0;
disk_mem[13877] = 0;
disk_mem[13878] = 0;
disk_mem[13879] = 0;
disk_mem[13880] = 0;
disk_mem[13881] = 0;
disk_mem[13882] = 0;
disk_mem[13883] = 0;
disk_mem[13884] = 0;
disk_mem[13885] = 0;
disk_mem[13886] = 0;
disk_mem[13887] = 0;
disk_mem[13888] = 0;
disk_mem[13889] = 0;
disk_mem[13890] = 0;
disk_mem[13891] = 0;
disk_mem[13892] = 0;
disk_mem[13893] = 0;
disk_mem[13894] = 0;
disk_mem[13895] = 0;
disk_mem[13896] = 0;
disk_mem[13897] = 0;
disk_mem[13898] = 0;
disk_mem[13899] = 0;
disk_mem[13900] = 0;
disk_mem[13901] = 0;
disk_mem[13902] = 0;
disk_mem[13903] = 0;
disk_mem[13904] = 0;
disk_mem[13905] = 0;
disk_mem[13906] = 0;
disk_mem[13907] = 0;
disk_mem[13908] = 0;
disk_mem[13909] = 0;
disk_mem[13910] = 0;
disk_mem[13911] = 0;
disk_mem[13912] = 0;
disk_mem[13913] = 0;
disk_mem[13914] = 0;
disk_mem[13915] = 0;
disk_mem[13916] = 0;
disk_mem[13917] = 0;
disk_mem[13918] = 0;
disk_mem[13919] = 0;
disk_mem[13920] = 0;
disk_mem[13921] = 0;
disk_mem[13922] = 0;
disk_mem[13923] = 0;
disk_mem[13924] = 0;
disk_mem[13925] = 0;
disk_mem[13926] = 0;
disk_mem[13927] = 0;
disk_mem[13928] = 0;
disk_mem[13929] = 0;
disk_mem[13930] = 0;
disk_mem[13931] = 0;
disk_mem[13932] = 0;
disk_mem[13933] = 0;
disk_mem[13934] = 0;
disk_mem[13935] = 0;
disk_mem[13936] = 0;
disk_mem[13937] = 0;
disk_mem[13938] = 0;
disk_mem[13939] = 0;
disk_mem[13940] = 0;
disk_mem[13941] = 0;
disk_mem[13942] = 0;
disk_mem[13943] = 0;
disk_mem[13944] = 0;
disk_mem[13945] = 0;
disk_mem[13946] = 0;
disk_mem[13947] = 0;
disk_mem[13948] = 0;
disk_mem[13949] = 0;
disk_mem[13950] = 0;
disk_mem[13951] = 0;
disk_mem[13952] = 0;
disk_mem[13953] = 0;
disk_mem[13954] = 0;
disk_mem[13955] = 0;
disk_mem[13956] = 0;
disk_mem[13957] = 0;
disk_mem[13958] = 0;
disk_mem[13959] = 0;
disk_mem[13960] = 0;
disk_mem[13961] = 0;
disk_mem[13962] = 0;
disk_mem[13963] = 0;
disk_mem[13964] = 0;
disk_mem[13965] = 0;
disk_mem[13966] = 0;
disk_mem[13967] = 0;
disk_mem[13968] = 0;
disk_mem[13969] = 0;
disk_mem[13970] = 0;
disk_mem[13971] = 0;
disk_mem[13972] = 0;
disk_mem[13973] = 0;
disk_mem[13974] = 0;
disk_mem[13975] = 0;
disk_mem[13976] = 0;
disk_mem[13977] = 0;
disk_mem[13978] = 0;
disk_mem[13979] = 0;
disk_mem[13980] = 0;
disk_mem[13981] = 0;
disk_mem[13982] = 0;
disk_mem[13983] = 0;
disk_mem[13984] = 0;
disk_mem[13985] = 0;
disk_mem[13986] = 0;
disk_mem[13987] = 0;
disk_mem[13988] = 0;
disk_mem[13989] = 0;
disk_mem[13990] = 0;
disk_mem[13991] = 0;
disk_mem[13992] = 0;
disk_mem[13993] = 0;
disk_mem[13994] = 0;
disk_mem[13995] = 0;
disk_mem[13996] = 0;
disk_mem[13997] = 0;
disk_mem[13998] = 0;
disk_mem[13999] = 0;
disk_mem[14000] = 0;
disk_mem[14001] = 0;
disk_mem[14002] = 0;
disk_mem[14003] = 0;
disk_mem[14004] = 0;
disk_mem[14005] = 0;
disk_mem[14006] = 0;
disk_mem[14007] = 0;
disk_mem[14008] = 0;
disk_mem[14009] = 0;
disk_mem[14010] = 0;
disk_mem[14011] = 0;
disk_mem[14012] = 0;
disk_mem[14013] = 0;
disk_mem[14014] = 0;
disk_mem[14015] = 0;
disk_mem[14016] = 0;
disk_mem[14017] = 0;
disk_mem[14018] = 0;
disk_mem[14019] = 0;
disk_mem[14020] = 0;
disk_mem[14021] = 0;
disk_mem[14022] = 0;
disk_mem[14023] = 0;
disk_mem[14024] = 0;
disk_mem[14025] = 0;
disk_mem[14026] = 0;
disk_mem[14027] = 0;
disk_mem[14028] = 0;
disk_mem[14029] = 0;
disk_mem[14030] = 0;
disk_mem[14031] = 0;
disk_mem[14032] = 0;
disk_mem[14033] = 0;
disk_mem[14034] = 0;
disk_mem[14035] = 0;
disk_mem[14036] = 0;
disk_mem[14037] = 0;
disk_mem[14038] = 0;
disk_mem[14039] = 0;
disk_mem[14040] = 0;
disk_mem[14041] = 0;
disk_mem[14042] = 0;
disk_mem[14043] = 0;
disk_mem[14044] = 0;
disk_mem[14045] = 0;
disk_mem[14046] = 0;
disk_mem[14047] = 0;
disk_mem[14048] = 0;
disk_mem[14049] = 0;
disk_mem[14050] = 0;
disk_mem[14051] = 0;
disk_mem[14052] = 0;
disk_mem[14053] = 0;
disk_mem[14054] = 0;
disk_mem[14055] = 0;
disk_mem[14056] = 0;
disk_mem[14057] = 0;
disk_mem[14058] = 0;
disk_mem[14059] = 0;
disk_mem[14060] = 0;
disk_mem[14061] = 0;
disk_mem[14062] = 0;
disk_mem[14063] = 0;
disk_mem[14064] = 0;
disk_mem[14065] = 0;
disk_mem[14066] = 0;
disk_mem[14067] = 0;
disk_mem[14068] = 0;
disk_mem[14069] = 0;
disk_mem[14070] = 0;
disk_mem[14071] = 0;
disk_mem[14072] = 0;
disk_mem[14073] = 0;
disk_mem[14074] = 0;
disk_mem[14075] = 0;
disk_mem[14076] = 0;
disk_mem[14077] = 0;
disk_mem[14078] = 0;
disk_mem[14079] = 0;
disk_mem[14080] = 0;
disk_mem[14081] = 0;
disk_mem[14082] = 0;
disk_mem[14083] = 0;
disk_mem[14084] = 0;
disk_mem[14085] = 0;
disk_mem[14086] = 0;
disk_mem[14087] = 0;
disk_mem[14088] = 0;
disk_mem[14089] = 0;
disk_mem[14090] = 0;
disk_mem[14091] = 0;
disk_mem[14092] = 0;
disk_mem[14093] = 0;
disk_mem[14094] = 0;
disk_mem[14095] = 0;
disk_mem[14096] = 0;
disk_mem[14097] = 0;
disk_mem[14098] = 0;
disk_mem[14099] = 0;
disk_mem[14100] = 0;
disk_mem[14101] = 0;
disk_mem[14102] = 0;
disk_mem[14103] = 0;
disk_mem[14104] = 0;
disk_mem[14105] = 0;
disk_mem[14106] = 0;
disk_mem[14107] = 0;
disk_mem[14108] = 0;
disk_mem[14109] = 0;
disk_mem[14110] = 0;
disk_mem[14111] = 0;
disk_mem[14112] = 0;
disk_mem[14113] = 0;
disk_mem[14114] = 0;
disk_mem[14115] = 0;
disk_mem[14116] = 0;
disk_mem[14117] = 0;
disk_mem[14118] = 0;
disk_mem[14119] = 0;
disk_mem[14120] = 0;
disk_mem[14121] = 0;
disk_mem[14122] = 0;
disk_mem[14123] = 0;
disk_mem[14124] = 0;
disk_mem[14125] = 0;
disk_mem[14126] = 0;
disk_mem[14127] = 0;
disk_mem[14128] = 0;
disk_mem[14129] = 0;
disk_mem[14130] = 0;
disk_mem[14131] = 0;
disk_mem[14132] = 0;
disk_mem[14133] = 0;
disk_mem[14134] = 0;
disk_mem[14135] = 0;
disk_mem[14136] = 0;
disk_mem[14137] = 0;
disk_mem[14138] = 0;
disk_mem[14139] = 0;
disk_mem[14140] = 0;
disk_mem[14141] = 0;
disk_mem[14142] = 0;
disk_mem[14143] = 0;
disk_mem[14144] = 0;
disk_mem[14145] = 0;
disk_mem[14146] = 0;
disk_mem[14147] = 0;
disk_mem[14148] = 0;
disk_mem[14149] = 0;
disk_mem[14150] = 0;
disk_mem[14151] = 0;
disk_mem[14152] = 0;
disk_mem[14153] = 0;
disk_mem[14154] = 0;
disk_mem[14155] = 0;
disk_mem[14156] = 0;
disk_mem[14157] = 0;
disk_mem[14158] = 0;
disk_mem[14159] = 0;
disk_mem[14160] = 0;
disk_mem[14161] = 0;
disk_mem[14162] = 0;
disk_mem[14163] = 0;
disk_mem[14164] = 0;
disk_mem[14165] = 0;
disk_mem[14166] = 0;
disk_mem[14167] = 0;
disk_mem[14168] = 0;
disk_mem[14169] = 0;
disk_mem[14170] = 0;
disk_mem[14171] = 0;
disk_mem[14172] = 0;
disk_mem[14173] = 0;
disk_mem[14174] = 0;
disk_mem[14175] = 0;
disk_mem[14176] = 0;
disk_mem[14177] = 0;
disk_mem[14178] = 0;
disk_mem[14179] = 0;
disk_mem[14180] = 0;
disk_mem[14181] = 0;
disk_mem[14182] = 0;
disk_mem[14183] = 0;
disk_mem[14184] = 0;
disk_mem[14185] = 0;
disk_mem[14186] = 0;
disk_mem[14187] = 0;
disk_mem[14188] = 0;
disk_mem[14189] = 0;
disk_mem[14190] = 0;
disk_mem[14191] = 0;
disk_mem[14192] = 0;
disk_mem[14193] = 0;
disk_mem[14194] = 0;
disk_mem[14195] = 0;
disk_mem[14196] = 0;
disk_mem[14197] = 0;
disk_mem[14198] = 0;
disk_mem[14199] = 0;
disk_mem[14200] = 0;
disk_mem[14201] = 0;
disk_mem[14202] = 0;
disk_mem[14203] = 0;
disk_mem[14204] = 0;
disk_mem[14205] = 0;
disk_mem[14206] = 0;
disk_mem[14207] = 0;
disk_mem[14208] = 0;
disk_mem[14209] = 0;
disk_mem[14210] = 0;
disk_mem[14211] = 0;
disk_mem[14212] = 0;
disk_mem[14213] = 0;
disk_mem[14214] = 0;
disk_mem[14215] = 0;
disk_mem[14216] = 0;
disk_mem[14217] = 0;
disk_mem[14218] = 0;
disk_mem[14219] = 0;
disk_mem[14220] = 0;
disk_mem[14221] = 0;
disk_mem[14222] = 0;
disk_mem[14223] = 0;
disk_mem[14224] = 0;
disk_mem[14225] = 0;
disk_mem[14226] = 0;
disk_mem[14227] = 0;
disk_mem[14228] = 0;
disk_mem[14229] = 0;
disk_mem[14230] = 0;
disk_mem[14231] = 0;
disk_mem[14232] = 0;
disk_mem[14233] = 0;
disk_mem[14234] = 0;
disk_mem[14235] = 0;
disk_mem[14236] = 0;
disk_mem[14237] = 0;
disk_mem[14238] = 0;
disk_mem[14239] = 0;
disk_mem[14240] = 0;
disk_mem[14241] = 0;
disk_mem[14242] = 0;
disk_mem[14243] = 0;
disk_mem[14244] = 0;
disk_mem[14245] = 0;
disk_mem[14246] = 0;
disk_mem[14247] = 0;
disk_mem[14248] = 0;
disk_mem[14249] = 0;
disk_mem[14250] = 0;
disk_mem[14251] = 0;
disk_mem[14252] = 0;
disk_mem[14253] = 0;
disk_mem[14254] = 0;
disk_mem[14255] = 0;
disk_mem[14256] = 0;
disk_mem[14257] = 0;
disk_mem[14258] = 0;
disk_mem[14259] = 0;
disk_mem[14260] = 0;
disk_mem[14261] = 0;
disk_mem[14262] = 0;
disk_mem[14263] = 0;
disk_mem[14264] = 0;
disk_mem[14265] = 0;
disk_mem[14266] = 0;
disk_mem[14267] = 0;
disk_mem[14268] = 0;
disk_mem[14269] = 0;
disk_mem[14270] = 0;
disk_mem[14271] = 0;
disk_mem[14272] = 0;
disk_mem[14273] = 0;
disk_mem[14274] = 0;
disk_mem[14275] = 0;
disk_mem[14276] = 0;
disk_mem[14277] = 0;
disk_mem[14278] = 0;
disk_mem[14279] = 0;
disk_mem[14280] = 0;
disk_mem[14281] = 0;
disk_mem[14282] = 0;
disk_mem[14283] = 0;
disk_mem[14284] = 0;
disk_mem[14285] = 0;
disk_mem[14286] = 0;
disk_mem[14287] = 0;
disk_mem[14288] = 0;
disk_mem[14289] = 0;
disk_mem[14290] = 0;
disk_mem[14291] = 0;
disk_mem[14292] = 0;
disk_mem[14293] = 0;
disk_mem[14294] = 0;
disk_mem[14295] = 0;
disk_mem[14296] = 0;
disk_mem[14297] = 0;
disk_mem[14298] = 0;
disk_mem[14299] = 0;
disk_mem[14300] = 0;
disk_mem[14301] = 0;
disk_mem[14302] = 0;
disk_mem[14303] = 0;
disk_mem[14304] = 0;
disk_mem[14305] = 0;
disk_mem[14306] = 0;
disk_mem[14307] = 0;
disk_mem[14308] = 0;
disk_mem[14309] = 0;
disk_mem[14310] = 0;
disk_mem[14311] = 0;
disk_mem[14312] = 0;
disk_mem[14313] = 0;
disk_mem[14314] = 0;
disk_mem[14315] = 0;
disk_mem[14316] = 0;
disk_mem[14317] = 0;
disk_mem[14318] = 0;
disk_mem[14319] = 0;
disk_mem[14320] = 0;
disk_mem[14321] = 0;
disk_mem[14322] = 0;
disk_mem[14323] = 0;
disk_mem[14324] = 0;
disk_mem[14325] = 0;
disk_mem[14326] = 0;
disk_mem[14327] = 0;
disk_mem[14328] = 0;
disk_mem[14329] = 0;
disk_mem[14330] = 0;
disk_mem[14331] = 0;
disk_mem[14332] = 0;
disk_mem[14333] = 0;
disk_mem[14334] = 0;
disk_mem[14335] = 0;
disk_mem[14336] = 0;
disk_mem[14337] = 0;
disk_mem[14338] = 0;
disk_mem[14339] = 0;
disk_mem[14340] = 0;
disk_mem[14341] = 0;
disk_mem[14342] = 0;
disk_mem[14343] = 0;
disk_mem[14344] = 0;
disk_mem[14345] = 0;
disk_mem[14346] = 0;
disk_mem[14347] = 0;
disk_mem[14348] = 0;
disk_mem[14349] = 0;
disk_mem[14350] = 0;
disk_mem[14351] = 0;
disk_mem[14352] = 0;
disk_mem[14353] = 0;
disk_mem[14354] = 0;
disk_mem[14355] = 0;
disk_mem[14356] = 0;
disk_mem[14357] = 0;
disk_mem[14358] = 0;
disk_mem[14359] = 0;
disk_mem[14360] = 0;
disk_mem[14361] = 0;
disk_mem[14362] = 0;
disk_mem[14363] = 0;
disk_mem[14364] = 0;
disk_mem[14365] = 0;
disk_mem[14366] = 0;
disk_mem[14367] = 0;
disk_mem[14368] = 0;
disk_mem[14369] = 0;
disk_mem[14370] = 0;
disk_mem[14371] = 0;
disk_mem[14372] = 0;
disk_mem[14373] = 0;
disk_mem[14374] = 0;
disk_mem[14375] = 0;
disk_mem[14376] = 0;
disk_mem[14377] = 0;
disk_mem[14378] = 0;
disk_mem[14379] = 0;
disk_mem[14380] = 0;
disk_mem[14381] = 0;
disk_mem[14382] = 0;
disk_mem[14383] = 0;
disk_mem[14384] = 0;
disk_mem[14385] = 0;
disk_mem[14386] = 0;
disk_mem[14387] = 0;
disk_mem[14388] = 0;
disk_mem[14389] = 0;
disk_mem[14390] = 0;
disk_mem[14391] = 0;
disk_mem[14392] = 0;
disk_mem[14393] = 0;
disk_mem[14394] = 0;
disk_mem[14395] = 0;
disk_mem[14396] = 0;
disk_mem[14397] = 0;
disk_mem[14398] = 0;
disk_mem[14399] = 0;
disk_mem[14400] = 0;
disk_mem[14401] = 0;
disk_mem[14402] = 0;
disk_mem[14403] = 0;
disk_mem[14404] = 0;
disk_mem[14405] = 0;
disk_mem[14406] = 0;
disk_mem[14407] = 0;
disk_mem[14408] = 0;
disk_mem[14409] = 0;
disk_mem[14410] = 0;
disk_mem[14411] = 0;
disk_mem[14412] = 0;
disk_mem[14413] = 0;
disk_mem[14414] = 0;
disk_mem[14415] = 0;
disk_mem[14416] = 0;
disk_mem[14417] = 0;
disk_mem[14418] = 0;
disk_mem[14419] = 0;
disk_mem[14420] = 0;
disk_mem[14421] = 0;
disk_mem[14422] = 0;
disk_mem[14423] = 0;
disk_mem[14424] = 0;
disk_mem[14425] = 0;
disk_mem[14426] = 0;
disk_mem[14427] = 0;
disk_mem[14428] = 0;
disk_mem[14429] = 0;
disk_mem[14430] = 0;
disk_mem[14431] = 0;
disk_mem[14432] = 0;
disk_mem[14433] = 0;
disk_mem[14434] = 0;
disk_mem[14435] = 0;
disk_mem[14436] = 0;
disk_mem[14437] = 0;
disk_mem[14438] = 0;
disk_mem[14439] = 0;
disk_mem[14440] = 0;
disk_mem[14441] = 0;
disk_mem[14442] = 0;
disk_mem[14443] = 0;
disk_mem[14444] = 0;
disk_mem[14445] = 0;
disk_mem[14446] = 0;
disk_mem[14447] = 0;
disk_mem[14448] = 0;
disk_mem[14449] = 0;
disk_mem[14450] = 0;
disk_mem[14451] = 0;
disk_mem[14452] = 0;
disk_mem[14453] = 0;
disk_mem[14454] = 0;
disk_mem[14455] = 0;
disk_mem[14456] = 0;
disk_mem[14457] = 0;
disk_mem[14458] = 0;
disk_mem[14459] = 0;
disk_mem[14460] = 0;
disk_mem[14461] = 0;
disk_mem[14462] = 0;
disk_mem[14463] = 0;
disk_mem[14464] = 0;
disk_mem[14465] = 0;
disk_mem[14466] = 0;
disk_mem[14467] = 0;
disk_mem[14468] = 0;
disk_mem[14469] = 0;
disk_mem[14470] = 0;
disk_mem[14471] = 0;
disk_mem[14472] = 0;
disk_mem[14473] = 0;
disk_mem[14474] = 0;
disk_mem[14475] = 0;
disk_mem[14476] = 0;
disk_mem[14477] = 0;
disk_mem[14478] = 0;
disk_mem[14479] = 0;
disk_mem[14480] = 0;
disk_mem[14481] = 0;
disk_mem[14482] = 0;
disk_mem[14483] = 0;
disk_mem[14484] = 0;
disk_mem[14485] = 0;
disk_mem[14486] = 0;
disk_mem[14487] = 0;
disk_mem[14488] = 0;
disk_mem[14489] = 0;
disk_mem[14490] = 0;
disk_mem[14491] = 0;
disk_mem[14492] = 0;
disk_mem[14493] = 0;
disk_mem[14494] = 0;
disk_mem[14495] = 0;
disk_mem[14496] = 0;
disk_mem[14497] = 0;
disk_mem[14498] = 0;
disk_mem[14499] = 0;
disk_mem[14500] = 0;
disk_mem[14501] = 0;
disk_mem[14502] = 0;
disk_mem[14503] = 0;
disk_mem[14504] = 0;
disk_mem[14505] = 0;
disk_mem[14506] = 0;
disk_mem[14507] = 0;
disk_mem[14508] = 0;
disk_mem[14509] = 0;
disk_mem[14510] = 0;
disk_mem[14511] = 0;
disk_mem[14512] = 0;
disk_mem[14513] = 0;
disk_mem[14514] = 0;
disk_mem[14515] = 0;
disk_mem[14516] = 0;
disk_mem[14517] = 0;
disk_mem[14518] = 0;
disk_mem[14519] = 0;
disk_mem[14520] = 0;
disk_mem[14521] = 0;
disk_mem[14522] = 0;
disk_mem[14523] = 0;
disk_mem[14524] = 0;
disk_mem[14525] = 0;
disk_mem[14526] = 0;
disk_mem[14527] = 0;
disk_mem[14528] = 0;
disk_mem[14529] = 0;
disk_mem[14530] = 0;
disk_mem[14531] = 0;
disk_mem[14532] = 0;
disk_mem[14533] = 0;
disk_mem[14534] = 0;
disk_mem[14535] = 0;
disk_mem[14536] = 0;
disk_mem[14537] = 0;
disk_mem[14538] = 0;
disk_mem[14539] = 0;
disk_mem[14540] = 0;
disk_mem[14541] = 0;
disk_mem[14542] = 0;
disk_mem[14543] = 0;
disk_mem[14544] = 0;
disk_mem[14545] = 0;
disk_mem[14546] = 0;
disk_mem[14547] = 0;
disk_mem[14548] = 0;
disk_mem[14549] = 0;
disk_mem[14550] = 0;
disk_mem[14551] = 0;
disk_mem[14552] = 0;
disk_mem[14553] = 0;
disk_mem[14554] = 0;
disk_mem[14555] = 0;
disk_mem[14556] = 0;
disk_mem[14557] = 0;
disk_mem[14558] = 0;
disk_mem[14559] = 0;
disk_mem[14560] = 0;
disk_mem[14561] = 0;
disk_mem[14562] = 0;
disk_mem[14563] = 0;
disk_mem[14564] = 0;
disk_mem[14565] = 0;
disk_mem[14566] = 0;
disk_mem[14567] = 0;
disk_mem[14568] = 0;
disk_mem[14569] = 0;
disk_mem[14570] = 0;
disk_mem[14571] = 0;
disk_mem[14572] = 0;
disk_mem[14573] = 0;
disk_mem[14574] = 0;
disk_mem[14575] = 0;
disk_mem[14576] = 0;
disk_mem[14577] = 0;
disk_mem[14578] = 0;
disk_mem[14579] = 0;
disk_mem[14580] = 0;
disk_mem[14581] = 0;
disk_mem[14582] = 0;
disk_mem[14583] = 0;
disk_mem[14584] = 0;
disk_mem[14585] = 0;
disk_mem[14586] = 0;
disk_mem[14587] = 0;
disk_mem[14588] = 0;
disk_mem[14589] = 0;
disk_mem[14590] = 0;
disk_mem[14591] = 0;
disk_mem[14592] = 0;
disk_mem[14593] = 0;
disk_mem[14594] = 0;
disk_mem[14595] = 0;
disk_mem[14596] = 0;
disk_mem[14597] = 0;
disk_mem[14598] = 0;
disk_mem[14599] = 0;
disk_mem[14600] = 0;
disk_mem[14601] = 0;
disk_mem[14602] = 0;
disk_mem[14603] = 0;
disk_mem[14604] = 0;
disk_mem[14605] = 0;
disk_mem[14606] = 0;
disk_mem[14607] = 0;
disk_mem[14608] = 0;
disk_mem[14609] = 0;
disk_mem[14610] = 0;
disk_mem[14611] = 0;
disk_mem[14612] = 0;
disk_mem[14613] = 0;
disk_mem[14614] = 0;
disk_mem[14615] = 0;
disk_mem[14616] = 0;
disk_mem[14617] = 0;
disk_mem[14618] = 0;
disk_mem[14619] = 0;
disk_mem[14620] = 0;
disk_mem[14621] = 0;
disk_mem[14622] = 0;
disk_mem[14623] = 0;
disk_mem[14624] = 0;
disk_mem[14625] = 0;
disk_mem[14626] = 0;
disk_mem[14627] = 0;
disk_mem[14628] = 0;
disk_mem[14629] = 0;
disk_mem[14630] = 0;
disk_mem[14631] = 0;
disk_mem[14632] = 0;
disk_mem[14633] = 0;
disk_mem[14634] = 0;
disk_mem[14635] = 0;
disk_mem[14636] = 0;
disk_mem[14637] = 0;
disk_mem[14638] = 0;
disk_mem[14639] = 0;
disk_mem[14640] = 0;
disk_mem[14641] = 0;
disk_mem[14642] = 0;
disk_mem[14643] = 0;
disk_mem[14644] = 0;
disk_mem[14645] = 0;
disk_mem[14646] = 0;
disk_mem[14647] = 0;
disk_mem[14648] = 0;
disk_mem[14649] = 0;
disk_mem[14650] = 0;
disk_mem[14651] = 0;
disk_mem[14652] = 0;
disk_mem[14653] = 0;
disk_mem[14654] = 0;
disk_mem[14655] = 0;
disk_mem[14656] = 0;
disk_mem[14657] = 0;
disk_mem[14658] = 0;
disk_mem[14659] = 0;
disk_mem[14660] = 0;
disk_mem[14661] = 0;
disk_mem[14662] = 0;
disk_mem[14663] = 0;
disk_mem[14664] = 0;
disk_mem[14665] = 0;
disk_mem[14666] = 0;
disk_mem[14667] = 0;
disk_mem[14668] = 0;
disk_mem[14669] = 0;
disk_mem[14670] = 0;
disk_mem[14671] = 0;
disk_mem[14672] = 0;
disk_mem[14673] = 0;
disk_mem[14674] = 0;
disk_mem[14675] = 0;
disk_mem[14676] = 0;
disk_mem[14677] = 0;
disk_mem[14678] = 0;
disk_mem[14679] = 0;
disk_mem[14680] = 0;
disk_mem[14681] = 0;
disk_mem[14682] = 0;
disk_mem[14683] = 0;
disk_mem[14684] = 0;
disk_mem[14685] = 0;
disk_mem[14686] = 0;
disk_mem[14687] = 0;
disk_mem[14688] = 0;
disk_mem[14689] = 0;
disk_mem[14690] = 0;
disk_mem[14691] = 0;
disk_mem[14692] = 0;
disk_mem[14693] = 0;
disk_mem[14694] = 0;
disk_mem[14695] = 0;
disk_mem[14696] = 0;
disk_mem[14697] = 0;
disk_mem[14698] = 0;
disk_mem[14699] = 0;
disk_mem[14700] = 0;
disk_mem[14701] = 0;
disk_mem[14702] = 0;
disk_mem[14703] = 0;
disk_mem[14704] = 0;
disk_mem[14705] = 0;
disk_mem[14706] = 0;
disk_mem[14707] = 0;
disk_mem[14708] = 0;
disk_mem[14709] = 0;
disk_mem[14710] = 0;
disk_mem[14711] = 0;
disk_mem[14712] = 0;
disk_mem[14713] = 0;
disk_mem[14714] = 0;
disk_mem[14715] = 0;
disk_mem[14716] = 0;
disk_mem[14717] = 0;
disk_mem[14718] = 0;
disk_mem[14719] = 0;
disk_mem[14720] = 0;
disk_mem[14721] = 0;
disk_mem[14722] = 0;
disk_mem[14723] = 0;
disk_mem[14724] = 0;
disk_mem[14725] = 0;
disk_mem[14726] = 0;
disk_mem[14727] = 0;
disk_mem[14728] = 0;
disk_mem[14729] = 0;
disk_mem[14730] = 0;
disk_mem[14731] = 0;
disk_mem[14732] = 0;
disk_mem[14733] = 0;
disk_mem[14734] = 0;
disk_mem[14735] = 0;
disk_mem[14736] = 0;
disk_mem[14737] = 0;
disk_mem[14738] = 0;
disk_mem[14739] = 0;
disk_mem[14740] = 0;
disk_mem[14741] = 0;
disk_mem[14742] = 0;
disk_mem[14743] = 0;
disk_mem[14744] = 0;
disk_mem[14745] = 0;
disk_mem[14746] = 0;
disk_mem[14747] = 0;
disk_mem[14748] = 0;
disk_mem[14749] = 0;
disk_mem[14750] = 0;
disk_mem[14751] = 0;
disk_mem[14752] = 0;
disk_mem[14753] = 0;
disk_mem[14754] = 0;
disk_mem[14755] = 0;
disk_mem[14756] = 0;
disk_mem[14757] = 0;
disk_mem[14758] = 0;
disk_mem[14759] = 0;
disk_mem[14760] = 0;
disk_mem[14761] = 0;
disk_mem[14762] = 0;
disk_mem[14763] = 0;
disk_mem[14764] = 0;
disk_mem[14765] = 0;
disk_mem[14766] = 0;
disk_mem[14767] = 0;
disk_mem[14768] = 0;
disk_mem[14769] = 0;
disk_mem[14770] = 0;
disk_mem[14771] = 0;
disk_mem[14772] = 0;
disk_mem[14773] = 0;
disk_mem[14774] = 0;
disk_mem[14775] = 0;
disk_mem[14776] = 0;
disk_mem[14777] = 0;
disk_mem[14778] = 0;
disk_mem[14779] = 0;
disk_mem[14780] = 0;
disk_mem[14781] = 0;
disk_mem[14782] = 0;
disk_mem[14783] = 0;
disk_mem[14784] = 0;
disk_mem[14785] = 0;
disk_mem[14786] = 0;
disk_mem[14787] = 0;
disk_mem[14788] = 0;
disk_mem[14789] = 0;
disk_mem[14790] = 0;
disk_mem[14791] = 0;
disk_mem[14792] = 0;
disk_mem[14793] = 0;
disk_mem[14794] = 0;
disk_mem[14795] = 0;
disk_mem[14796] = 0;
disk_mem[14797] = 0;
disk_mem[14798] = 0;
disk_mem[14799] = 0;
disk_mem[14800] = 0;
disk_mem[14801] = 0;
disk_mem[14802] = 0;
disk_mem[14803] = 0;
disk_mem[14804] = 0;
disk_mem[14805] = 0;
disk_mem[14806] = 0;
disk_mem[14807] = 0;
disk_mem[14808] = 0;
disk_mem[14809] = 0;
disk_mem[14810] = 0;
disk_mem[14811] = 0;
disk_mem[14812] = 0;
disk_mem[14813] = 0;
disk_mem[14814] = 0;
disk_mem[14815] = 0;
disk_mem[14816] = 0;
disk_mem[14817] = 0;
disk_mem[14818] = 0;
disk_mem[14819] = 0;
disk_mem[14820] = 0;
disk_mem[14821] = 0;
disk_mem[14822] = 0;
disk_mem[14823] = 0;
disk_mem[14824] = 0;
disk_mem[14825] = 0;
disk_mem[14826] = 0;
disk_mem[14827] = 0;
disk_mem[14828] = 0;
disk_mem[14829] = 0;
disk_mem[14830] = 0;
disk_mem[14831] = 0;
disk_mem[14832] = 0;
disk_mem[14833] = 0;
disk_mem[14834] = 0;
disk_mem[14835] = 0;
disk_mem[14836] = 0;
disk_mem[14837] = 0;
disk_mem[14838] = 0;
disk_mem[14839] = 0;
disk_mem[14840] = 0;
disk_mem[14841] = 0;
disk_mem[14842] = 0;
disk_mem[14843] = 0;
disk_mem[14844] = 0;
disk_mem[14845] = 0;
disk_mem[14846] = 0;
disk_mem[14847] = 0;
disk_mem[14848] = 0;
disk_mem[14849] = 0;
disk_mem[14850] = 0;
disk_mem[14851] = 0;
disk_mem[14852] = 0;
disk_mem[14853] = 0;
disk_mem[14854] = 0;
disk_mem[14855] = 0;
disk_mem[14856] = 0;
disk_mem[14857] = 0;
disk_mem[14858] = 0;
disk_mem[14859] = 0;
disk_mem[14860] = 0;
disk_mem[14861] = 0;
disk_mem[14862] = 0;
disk_mem[14863] = 0;
disk_mem[14864] = 0;
disk_mem[14865] = 0;
disk_mem[14866] = 0;
disk_mem[14867] = 0;
disk_mem[14868] = 0;
disk_mem[14869] = 0;
disk_mem[14870] = 0;
disk_mem[14871] = 0;
disk_mem[14872] = 0;
disk_mem[14873] = 0;
disk_mem[14874] = 0;
disk_mem[14875] = 0;
disk_mem[14876] = 0;
disk_mem[14877] = 0;
disk_mem[14878] = 0;
disk_mem[14879] = 0;
disk_mem[14880] = 0;
disk_mem[14881] = 0;
disk_mem[14882] = 0;
disk_mem[14883] = 0;
disk_mem[14884] = 0;
disk_mem[14885] = 0;
disk_mem[14886] = 0;
disk_mem[14887] = 0;
disk_mem[14888] = 0;
disk_mem[14889] = 0;
disk_mem[14890] = 0;
disk_mem[14891] = 0;
disk_mem[14892] = 0;
disk_mem[14893] = 0;
disk_mem[14894] = 0;
disk_mem[14895] = 0;
disk_mem[14896] = 0;
disk_mem[14897] = 0;
disk_mem[14898] = 0;
disk_mem[14899] = 0;
disk_mem[14900] = 0;
disk_mem[14901] = 0;
disk_mem[14902] = 0;
disk_mem[14903] = 0;
disk_mem[14904] = 0;
disk_mem[14905] = 0;
disk_mem[14906] = 0;
disk_mem[14907] = 0;
disk_mem[14908] = 0;
disk_mem[14909] = 0;
disk_mem[14910] = 0;
disk_mem[14911] = 0;
disk_mem[14912] = 0;
disk_mem[14913] = 0;
disk_mem[14914] = 0;
disk_mem[14915] = 0;
disk_mem[14916] = 0;
disk_mem[14917] = 0;
disk_mem[14918] = 0;
disk_mem[14919] = 0;
disk_mem[14920] = 0;
disk_mem[14921] = 0;
disk_mem[14922] = 0;
disk_mem[14923] = 0;
disk_mem[14924] = 0;
disk_mem[14925] = 0;
disk_mem[14926] = 0;
disk_mem[14927] = 0;
disk_mem[14928] = 0;
disk_mem[14929] = 0;
disk_mem[14930] = 0;
disk_mem[14931] = 0;
disk_mem[14932] = 0;
disk_mem[14933] = 0;
disk_mem[14934] = 0;
disk_mem[14935] = 0;
disk_mem[14936] = 0;
disk_mem[14937] = 0;
disk_mem[14938] = 0;
disk_mem[14939] = 0;
disk_mem[14940] = 0;
disk_mem[14941] = 0;
disk_mem[14942] = 0;
disk_mem[14943] = 0;
disk_mem[14944] = 0;
disk_mem[14945] = 0;
disk_mem[14946] = 0;
disk_mem[14947] = 0;
disk_mem[14948] = 0;
disk_mem[14949] = 0;
disk_mem[14950] = 0;
disk_mem[14951] = 0;
disk_mem[14952] = 0;
disk_mem[14953] = 0;
disk_mem[14954] = 0;
disk_mem[14955] = 0;
disk_mem[14956] = 0;
disk_mem[14957] = 0;
disk_mem[14958] = 0;
disk_mem[14959] = 0;
disk_mem[14960] = 0;
disk_mem[14961] = 0;
disk_mem[14962] = 0;
disk_mem[14963] = 0;
disk_mem[14964] = 0;
disk_mem[14965] = 0;
disk_mem[14966] = 0;
disk_mem[14967] = 0;
disk_mem[14968] = 0;
disk_mem[14969] = 0;
disk_mem[14970] = 0;
disk_mem[14971] = 0;
disk_mem[14972] = 0;
disk_mem[14973] = 0;
disk_mem[14974] = 0;
disk_mem[14975] = 0;
disk_mem[14976] = 0;
disk_mem[14977] = 0;
disk_mem[14978] = 0;
disk_mem[14979] = 0;
disk_mem[14980] = 0;
disk_mem[14981] = 0;
disk_mem[14982] = 0;
disk_mem[14983] = 0;
disk_mem[14984] = 0;
disk_mem[14985] = 0;
disk_mem[14986] = 0;
disk_mem[14987] = 0;
disk_mem[14988] = 0;
disk_mem[14989] = 0;
disk_mem[14990] = 0;
disk_mem[14991] = 0;
disk_mem[14992] = 0;
disk_mem[14993] = 0;
disk_mem[14994] = 0;
disk_mem[14995] = 0;
disk_mem[14996] = 0;
disk_mem[14997] = 0;
disk_mem[14998] = 0;
disk_mem[14999] = 0;
disk_mem[15000] = 0;
disk_mem[15001] = 0;
disk_mem[15002] = 0;
disk_mem[15003] = 0;
disk_mem[15004] = 0;
disk_mem[15005] = 0;
disk_mem[15006] = 0;
disk_mem[15007] = 0;
disk_mem[15008] = 0;
disk_mem[15009] = 0;
disk_mem[15010] = 0;
disk_mem[15011] = 0;
disk_mem[15012] = 0;
disk_mem[15013] = 0;
disk_mem[15014] = 0;
disk_mem[15015] = 0;
disk_mem[15016] = 0;
disk_mem[15017] = 0;
disk_mem[15018] = 0;
disk_mem[15019] = 0;
disk_mem[15020] = 0;
disk_mem[15021] = 0;
disk_mem[15022] = 0;
disk_mem[15023] = 0;
disk_mem[15024] = 0;
disk_mem[15025] = 0;
disk_mem[15026] = 0;
disk_mem[15027] = 0;
disk_mem[15028] = 0;
disk_mem[15029] = 0;
disk_mem[15030] = 0;
disk_mem[15031] = 0;
disk_mem[15032] = 0;
disk_mem[15033] = 0;
disk_mem[15034] = 0;
disk_mem[15035] = 0;
disk_mem[15036] = 0;
disk_mem[15037] = 0;
disk_mem[15038] = 0;
disk_mem[15039] = 0;
disk_mem[15040] = 0;
disk_mem[15041] = 0;
disk_mem[15042] = 0;
disk_mem[15043] = 0;
disk_mem[15044] = 0;
disk_mem[15045] = 0;
disk_mem[15046] = 0;
disk_mem[15047] = 0;
disk_mem[15048] = 0;
disk_mem[15049] = 0;
disk_mem[15050] = 0;
disk_mem[15051] = 0;
disk_mem[15052] = 0;
disk_mem[15053] = 0;
disk_mem[15054] = 0;
disk_mem[15055] = 0;
disk_mem[15056] = 0;
disk_mem[15057] = 0;
disk_mem[15058] = 0;
disk_mem[15059] = 0;
disk_mem[15060] = 0;
disk_mem[15061] = 0;
disk_mem[15062] = 0;
disk_mem[15063] = 0;
disk_mem[15064] = 0;
disk_mem[15065] = 0;
disk_mem[15066] = 0;
disk_mem[15067] = 0;
disk_mem[15068] = 0;
disk_mem[15069] = 0;
disk_mem[15070] = 0;
disk_mem[15071] = 0;
disk_mem[15072] = 0;
disk_mem[15073] = 0;
disk_mem[15074] = 0;
disk_mem[15075] = 0;
disk_mem[15076] = 0;
disk_mem[15077] = 0;
disk_mem[15078] = 0;
disk_mem[15079] = 0;
disk_mem[15080] = 0;
disk_mem[15081] = 0;
disk_mem[15082] = 0;
disk_mem[15083] = 0;
disk_mem[15084] = 0;
disk_mem[15085] = 0;
disk_mem[15086] = 0;
disk_mem[15087] = 0;
disk_mem[15088] = 0;
disk_mem[15089] = 0;
disk_mem[15090] = 0;
disk_mem[15091] = 0;
disk_mem[15092] = 0;
disk_mem[15093] = 0;
disk_mem[15094] = 0;
disk_mem[15095] = 0;
disk_mem[15096] = 0;
disk_mem[15097] = 0;
disk_mem[15098] = 0;
disk_mem[15099] = 0;
disk_mem[15100] = 0;
disk_mem[15101] = 0;
disk_mem[15102] = 0;
disk_mem[15103] = 0;
disk_mem[15104] = 0;
disk_mem[15105] = 0;
disk_mem[15106] = 0;
disk_mem[15107] = 0;
disk_mem[15108] = 0;
disk_mem[15109] = 0;
disk_mem[15110] = 0;
disk_mem[15111] = 0;
disk_mem[15112] = 0;
disk_mem[15113] = 0;
disk_mem[15114] = 0;
disk_mem[15115] = 0;
disk_mem[15116] = 0;
disk_mem[15117] = 0;
disk_mem[15118] = 0;
disk_mem[15119] = 0;
disk_mem[15120] = 0;
disk_mem[15121] = 0;
disk_mem[15122] = 0;
disk_mem[15123] = 0;
disk_mem[15124] = 0;
disk_mem[15125] = 0;
disk_mem[15126] = 0;
disk_mem[15127] = 0;
disk_mem[15128] = 0;
disk_mem[15129] = 0;
disk_mem[15130] = 0;
disk_mem[15131] = 0;
disk_mem[15132] = 0;
disk_mem[15133] = 0;
disk_mem[15134] = 0;
disk_mem[15135] = 0;
disk_mem[15136] = 0;
disk_mem[15137] = 0;
disk_mem[15138] = 0;
disk_mem[15139] = 0;
disk_mem[15140] = 0;
disk_mem[15141] = 0;
disk_mem[15142] = 0;
disk_mem[15143] = 0;
disk_mem[15144] = 0;
disk_mem[15145] = 0;
disk_mem[15146] = 0;
disk_mem[15147] = 0;
disk_mem[15148] = 0;
disk_mem[15149] = 0;
disk_mem[15150] = 0;
disk_mem[15151] = 0;
disk_mem[15152] = 0;
disk_mem[15153] = 0;
disk_mem[15154] = 0;
disk_mem[15155] = 0;
disk_mem[15156] = 0;
disk_mem[15157] = 0;
disk_mem[15158] = 0;
disk_mem[15159] = 0;
disk_mem[15160] = 0;
disk_mem[15161] = 0;
disk_mem[15162] = 0;
disk_mem[15163] = 0;
disk_mem[15164] = 0;
disk_mem[15165] = 0;
disk_mem[15166] = 0;
disk_mem[15167] = 0;
disk_mem[15168] = 0;
disk_mem[15169] = 0;
disk_mem[15170] = 0;
disk_mem[15171] = 0;
disk_mem[15172] = 0;
disk_mem[15173] = 0;
disk_mem[15174] = 0;
disk_mem[15175] = 0;
disk_mem[15176] = 0;
disk_mem[15177] = 0;
disk_mem[15178] = 0;
disk_mem[15179] = 0;
disk_mem[15180] = 0;
disk_mem[15181] = 0;
disk_mem[15182] = 0;
disk_mem[15183] = 0;
disk_mem[15184] = 0;
disk_mem[15185] = 0;
disk_mem[15186] = 0;
disk_mem[15187] = 0;
disk_mem[15188] = 0;
disk_mem[15189] = 0;
disk_mem[15190] = 0;
disk_mem[15191] = 0;
disk_mem[15192] = 0;
disk_mem[15193] = 0;
disk_mem[15194] = 0;
disk_mem[15195] = 0;
disk_mem[15196] = 0;
disk_mem[15197] = 0;
disk_mem[15198] = 0;
disk_mem[15199] = 0;
disk_mem[15200] = 0;
disk_mem[15201] = 0;
disk_mem[15202] = 0;
disk_mem[15203] = 0;
disk_mem[15204] = 0;
disk_mem[15205] = 0;
disk_mem[15206] = 0;
disk_mem[15207] = 0;
disk_mem[15208] = 0;
disk_mem[15209] = 0;
disk_mem[15210] = 0;
disk_mem[15211] = 0;
disk_mem[15212] = 0;
disk_mem[15213] = 0;
disk_mem[15214] = 0;
disk_mem[15215] = 0;
disk_mem[15216] = 0;
disk_mem[15217] = 0;
disk_mem[15218] = 0;
disk_mem[15219] = 0;
disk_mem[15220] = 0;
disk_mem[15221] = 0;
disk_mem[15222] = 0;
disk_mem[15223] = 0;
disk_mem[15224] = 0;
disk_mem[15225] = 0;
disk_mem[15226] = 0;
disk_mem[15227] = 0;
disk_mem[15228] = 0;
disk_mem[15229] = 0;
disk_mem[15230] = 0;
disk_mem[15231] = 0;
disk_mem[15232] = 0;
disk_mem[15233] = 0;
disk_mem[15234] = 0;
disk_mem[15235] = 0;
disk_mem[15236] = 0;
disk_mem[15237] = 0;
disk_mem[15238] = 0;
disk_mem[15239] = 0;
disk_mem[15240] = 0;
disk_mem[15241] = 0;
disk_mem[15242] = 0;
disk_mem[15243] = 0;
disk_mem[15244] = 0;
disk_mem[15245] = 0;
disk_mem[15246] = 0;
disk_mem[15247] = 0;
disk_mem[15248] = 0;
disk_mem[15249] = 0;
disk_mem[15250] = 0;
disk_mem[15251] = 0;
disk_mem[15252] = 0;
disk_mem[15253] = 0;
disk_mem[15254] = 0;
disk_mem[15255] = 0;
disk_mem[15256] = 0;
disk_mem[15257] = 0;
disk_mem[15258] = 0;
disk_mem[15259] = 0;
disk_mem[15260] = 0;
disk_mem[15261] = 0;
disk_mem[15262] = 0;
disk_mem[15263] = 0;
disk_mem[15264] = 0;
disk_mem[15265] = 0;
disk_mem[15266] = 0;
disk_mem[15267] = 0;
disk_mem[15268] = 0;
disk_mem[15269] = 0;
disk_mem[15270] = 0;
disk_mem[15271] = 0;
disk_mem[15272] = 0;
disk_mem[15273] = 0;
disk_mem[15274] = 0;
disk_mem[15275] = 0;
disk_mem[15276] = 0;
disk_mem[15277] = 0;
disk_mem[15278] = 0;
disk_mem[15279] = 0;
disk_mem[15280] = 0;
disk_mem[15281] = 0;
disk_mem[15282] = 0;
disk_mem[15283] = 0;
disk_mem[15284] = 0;
disk_mem[15285] = 0;
disk_mem[15286] = 0;
disk_mem[15287] = 0;
disk_mem[15288] = 0;
disk_mem[15289] = 0;
disk_mem[15290] = 0;
disk_mem[15291] = 0;
disk_mem[15292] = 0;
disk_mem[15293] = 0;
disk_mem[15294] = 0;
disk_mem[15295] = 0;
disk_mem[15296] = 0;
disk_mem[15297] = 0;
disk_mem[15298] = 0;
disk_mem[15299] = 0;
disk_mem[15300] = 0;
disk_mem[15301] = 0;
disk_mem[15302] = 0;
disk_mem[15303] = 0;
disk_mem[15304] = 0;
disk_mem[15305] = 0;
disk_mem[15306] = 0;
disk_mem[15307] = 0;
disk_mem[15308] = 0;
disk_mem[15309] = 0;
disk_mem[15310] = 0;
disk_mem[15311] = 0;
disk_mem[15312] = 0;
disk_mem[15313] = 0;
disk_mem[15314] = 0;
disk_mem[15315] = 0;
disk_mem[15316] = 0;
disk_mem[15317] = 0;
disk_mem[15318] = 0;
disk_mem[15319] = 0;
disk_mem[15320] = 0;
disk_mem[15321] = 0;
disk_mem[15322] = 0;
disk_mem[15323] = 0;
disk_mem[15324] = 0;
disk_mem[15325] = 0;
disk_mem[15326] = 0;
disk_mem[15327] = 0;
disk_mem[15328] = 0;
disk_mem[15329] = 0;
disk_mem[15330] = 0;
disk_mem[15331] = 0;
disk_mem[15332] = 0;
disk_mem[15333] = 0;
disk_mem[15334] = 0;
disk_mem[15335] = 0;
disk_mem[15336] = 0;
disk_mem[15337] = 0;
disk_mem[15338] = 0;
disk_mem[15339] = 0;
disk_mem[15340] = 0;
disk_mem[15341] = 0;
disk_mem[15342] = 0;
disk_mem[15343] = 0;
disk_mem[15344] = 0;
disk_mem[15345] = 0;
disk_mem[15346] = 0;
disk_mem[15347] = 0;
disk_mem[15348] = 0;
disk_mem[15349] = 0;
disk_mem[15350] = 0;
disk_mem[15351] = 0;
disk_mem[15352] = 0;
disk_mem[15353] = 0;
disk_mem[15354] = 0;
disk_mem[15355] = 0;
disk_mem[15356] = 0;
disk_mem[15357] = 0;
disk_mem[15358] = 0;
disk_mem[15359] = 0;
disk_mem[15360] = 0;
disk_mem[15361] = 0;
disk_mem[15362] = 0;
disk_mem[15363] = 0;
disk_mem[15364] = 0;
disk_mem[15365] = 0;
disk_mem[15366] = 0;
disk_mem[15367] = 0;
disk_mem[15368] = 0;
disk_mem[15369] = 0;
disk_mem[15370] = 0;
disk_mem[15371] = 0;
disk_mem[15372] = 0;
disk_mem[15373] = 0;
disk_mem[15374] = 0;
disk_mem[15375] = 0;
disk_mem[15376] = 0;
disk_mem[15377] = 0;
disk_mem[15378] = 0;
disk_mem[15379] = 0;
disk_mem[15380] = 0;
disk_mem[15381] = 0;
disk_mem[15382] = 0;
disk_mem[15383] = 0;
disk_mem[15384] = 0;
disk_mem[15385] = 0;
disk_mem[15386] = 0;
disk_mem[15387] = 0;
disk_mem[15388] = 0;
disk_mem[15389] = 0;
disk_mem[15390] = 0;
disk_mem[15391] = 0;
disk_mem[15392] = 0;
disk_mem[15393] = 0;
disk_mem[15394] = 0;
disk_mem[15395] = 0;
disk_mem[15396] = 0;
disk_mem[15397] = 0;
disk_mem[15398] = 0;
disk_mem[15399] = 0;
disk_mem[15400] = 0;
disk_mem[15401] = 0;
disk_mem[15402] = 0;
disk_mem[15403] = 0;
disk_mem[15404] = 0;
disk_mem[15405] = 0;
disk_mem[15406] = 0;
disk_mem[15407] = 0;
disk_mem[15408] = 0;
disk_mem[15409] = 0;
disk_mem[15410] = 0;
disk_mem[15411] = 0;
disk_mem[15412] = 0;
disk_mem[15413] = 0;
disk_mem[15414] = 0;
disk_mem[15415] = 0;
disk_mem[15416] = 0;
disk_mem[15417] = 0;
disk_mem[15418] = 0;
disk_mem[15419] = 0;
disk_mem[15420] = 0;
disk_mem[15421] = 0;
disk_mem[15422] = 0;
disk_mem[15423] = 0;
disk_mem[15424] = 0;
disk_mem[15425] = 0;
disk_mem[15426] = 0;
disk_mem[15427] = 0;
disk_mem[15428] = 0;
disk_mem[15429] = 0;
disk_mem[15430] = 0;
disk_mem[15431] = 0;
disk_mem[15432] = 0;
disk_mem[15433] = 0;
disk_mem[15434] = 0;
disk_mem[15435] = 0;
disk_mem[15436] = 0;
disk_mem[15437] = 0;
disk_mem[15438] = 0;
disk_mem[15439] = 0;
disk_mem[15440] = 0;
disk_mem[15441] = 0;
disk_mem[15442] = 0;
disk_mem[15443] = 0;
disk_mem[15444] = 0;
disk_mem[15445] = 0;
disk_mem[15446] = 0;
disk_mem[15447] = 0;
disk_mem[15448] = 0;
disk_mem[15449] = 0;
disk_mem[15450] = 0;
disk_mem[15451] = 0;
disk_mem[15452] = 0;
disk_mem[15453] = 0;
disk_mem[15454] = 0;
disk_mem[15455] = 0;
disk_mem[15456] = 0;
disk_mem[15457] = 0;
disk_mem[15458] = 0;
disk_mem[15459] = 0;
disk_mem[15460] = 0;
disk_mem[15461] = 0;
disk_mem[15462] = 0;
disk_mem[15463] = 0;
disk_mem[15464] = 0;
disk_mem[15465] = 0;
disk_mem[15466] = 0;
disk_mem[15467] = 0;
disk_mem[15468] = 0;
disk_mem[15469] = 0;
disk_mem[15470] = 0;
disk_mem[15471] = 0;
disk_mem[15472] = 0;
disk_mem[15473] = 0;
disk_mem[15474] = 0;
disk_mem[15475] = 0;
disk_mem[15476] = 0;
disk_mem[15477] = 0;
disk_mem[15478] = 0;
disk_mem[15479] = 0;
disk_mem[15480] = 0;
disk_mem[15481] = 0;
disk_mem[15482] = 0;
disk_mem[15483] = 0;
disk_mem[15484] = 0;
disk_mem[15485] = 0;
disk_mem[15486] = 0;
disk_mem[15487] = 0;
disk_mem[15488] = 0;
disk_mem[15489] = 0;
disk_mem[15490] = 0;
disk_mem[15491] = 0;
disk_mem[15492] = 0;
disk_mem[15493] = 0;
disk_mem[15494] = 0;
disk_mem[15495] = 0;
disk_mem[15496] = 0;
disk_mem[15497] = 0;
disk_mem[15498] = 0;
disk_mem[15499] = 0;
disk_mem[15500] = 0;
disk_mem[15501] = 0;
disk_mem[15502] = 0;
disk_mem[15503] = 0;
disk_mem[15504] = 0;
disk_mem[15505] = 0;
disk_mem[15506] = 0;
disk_mem[15507] = 0;
disk_mem[15508] = 0;
disk_mem[15509] = 0;
disk_mem[15510] = 0;
disk_mem[15511] = 0;
disk_mem[15512] = 0;
disk_mem[15513] = 0;
disk_mem[15514] = 0;
disk_mem[15515] = 0;
disk_mem[15516] = 0;
disk_mem[15517] = 0;
disk_mem[15518] = 0;
disk_mem[15519] = 0;
disk_mem[15520] = 0;
disk_mem[15521] = 0;
disk_mem[15522] = 0;
disk_mem[15523] = 0;
disk_mem[15524] = 0;
disk_mem[15525] = 0;
disk_mem[15526] = 0;
disk_mem[15527] = 0;
disk_mem[15528] = 0;
disk_mem[15529] = 0;
disk_mem[15530] = 0;
disk_mem[15531] = 0;
disk_mem[15532] = 0;
disk_mem[15533] = 0;
disk_mem[15534] = 0;
disk_mem[15535] = 0;
disk_mem[15536] = 0;
disk_mem[15537] = 0;
disk_mem[15538] = 0;
disk_mem[15539] = 0;
disk_mem[15540] = 0;
disk_mem[15541] = 0;
disk_mem[15542] = 0;
disk_mem[15543] = 0;
disk_mem[15544] = 0;
disk_mem[15545] = 0;
disk_mem[15546] = 0;
disk_mem[15547] = 0;
disk_mem[15548] = 0;
disk_mem[15549] = 0;
disk_mem[15550] = 0;
disk_mem[15551] = 0;
disk_mem[15552] = 0;
disk_mem[15553] = 0;
disk_mem[15554] = 0;
disk_mem[15555] = 0;
disk_mem[15556] = 0;
disk_mem[15557] = 0;
disk_mem[15558] = 0;
disk_mem[15559] = 0;
disk_mem[15560] = 0;
disk_mem[15561] = 0;
disk_mem[15562] = 0;
disk_mem[15563] = 0;
disk_mem[15564] = 0;
disk_mem[15565] = 0;
disk_mem[15566] = 0;
disk_mem[15567] = 0;
disk_mem[15568] = 0;
disk_mem[15569] = 0;
disk_mem[15570] = 0;
disk_mem[15571] = 0;
disk_mem[15572] = 0;
disk_mem[15573] = 0;
disk_mem[15574] = 0;
disk_mem[15575] = 0;
disk_mem[15576] = 0;
disk_mem[15577] = 0;
disk_mem[15578] = 0;
disk_mem[15579] = 0;
disk_mem[15580] = 0;
disk_mem[15581] = 0;
disk_mem[15582] = 0;
disk_mem[15583] = 0;
disk_mem[15584] = 0;
disk_mem[15585] = 0;
disk_mem[15586] = 0;
disk_mem[15587] = 0;
disk_mem[15588] = 0;
disk_mem[15589] = 0;
disk_mem[15590] = 0;
disk_mem[15591] = 0;
disk_mem[15592] = 0;
disk_mem[15593] = 0;
disk_mem[15594] = 0;
disk_mem[15595] = 0;
disk_mem[15596] = 0;
disk_mem[15597] = 0;
disk_mem[15598] = 0;
disk_mem[15599] = 0;
disk_mem[15600] = 0;
disk_mem[15601] = 0;
disk_mem[15602] = 0;
disk_mem[15603] = 0;
disk_mem[15604] = 0;
disk_mem[15605] = 0;
disk_mem[15606] = 0;
disk_mem[15607] = 0;
disk_mem[15608] = 0;
disk_mem[15609] = 0;
disk_mem[15610] = 0;
disk_mem[15611] = 0;
disk_mem[15612] = 0;
disk_mem[15613] = 0;
disk_mem[15614] = 0;
disk_mem[15615] = 0;
disk_mem[15616] = 0;
disk_mem[15617] = 0;
disk_mem[15618] = 0;
disk_mem[15619] = 0;
disk_mem[15620] = 0;
disk_mem[15621] = 0;
disk_mem[15622] = 0;
disk_mem[15623] = 0;
disk_mem[15624] = 0;
disk_mem[15625] = 0;
disk_mem[15626] = 0;
disk_mem[15627] = 0;
disk_mem[15628] = 0;
disk_mem[15629] = 0;
disk_mem[15630] = 0;
disk_mem[15631] = 0;
disk_mem[15632] = 0;
disk_mem[15633] = 0;
disk_mem[15634] = 0;
disk_mem[15635] = 0;
disk_mem[15636] = 0;
disk_mem[15637] = 0;
disk_mem[15638] = 0;
disk_mem[15639] = 0;
disk_mem[15640] = 0;
disk_mem[15641] = 0;
disk_mem[15642] = 0;
disk_mem[15643] = 0;
disk_mem[15644] = 0;
disk_mem[15645] = 0;
disk_mem[15646] = 0;
disk_mem[15647] = 0;
disk_mem[15648] = 0;
disk_mem[15649] = 0;
disk_mem[15650] = 0;
disk_mem[15651] = 0;
disk_mem[15652] = 0;
disk_mem[15653] = 0;
disk_mem[15654] = 0;
disk_mem[15655] = 0;
disk_mem[15656] = 0;
disk_mem[15657] = 0;
disk_mem[15658] = 0;
disk_mem[15659] = 0;
disk_mem[15660] = 0;
disk_mem[15661] = 0;
disk_mem[15662] = 0;
disk_mem[15663] = 0;
disk_mem[15664] = 0;
disk_mem[15665] = 0;
disk_mem[15666] = 0;
disk_mem[15667] = 0;
disk_mem[15668] = 0;
disk_mem[15669] = 0;
disk_mem[15670] = 0;
disk_mem[15671] = 0;
disk_mem[15672] = 0;
disk_mem[15673] = 0;
disk_mem[15674] = 0;
disk_mem[15675] = 0;
disk_mem[15676] = 0;
disk_mem[15677] = 0;
disk_mem[15678] = 0;
disk_mem[15679] = 0;
disk_mem[15680] = 0;
disk_mem[15681] = 0;
disk_mem[15682] = 0;
disk_mem[15683] = 0;
disk_mem[15684] = 0;
disk_mem[15685] = 0;
disk_mem[15686] = 0;
disk_mem[15687] = 0;
disk_mem[15688] = 0;
disk_mem[15689] = 0;
disk_mem[15690] = 0;
disk_mem[15691] = 0;
disk_mem[15692] = 0;
disk_mem[15693] = 0;
disk_mem[15694] = 0;
disk_mem[15695] = 0;
disk_mem[15696] = 0;
disk_mem[15697] = 0;
disk_mem[15698] = 0;
disk_mem[15699] = 0;
disk_mem[15700] = 0;
disk_mem[15701] = 0;
disk_mem[15702] = 0;
disk_mem[15703] = 0;
disk_mem[15704] = 0;
disk_mem[15705] = 0;
disk_mem[15706] = 0;
disk_mem[15707] = 0;
disk_mem[15708] = 0;
disk_mem[15709] = 0;
disk_mem[15710] = 0;
disk_mem[15711] = 0;
disk_mem[15712] = 0;
disk_mem[15713] = 0;
disk_mem[15714] = 0;
disk_mem[15715] = 0;
disk_mem[15716] = 0;
disk_mem[15717] = 0;
disk_mem[15718] = 0;
disk_mem[15719] = 0;
disk_mem[15720] = 0;
disk_mem[15721] = 0;
disk_mem[15722] = 0;
disk_mem[15723] = 0;
disk_mem[15724] = 0;
disk_mem[15725] = 0;
disk_mem[15726] = 0;
disk_mem[15727] = 0;
disk_mem[15728] = 0;
disk_mem[15729] = 0;
disk_mem[15730] = 0;
disk_mem[15731] = 0;
disk_mem[15732] = 0;
disk_mem[15733] = 0;
disk_mem[15734] = 0;
disk_mem[15735] = 0;
disk_mem[15736] = 0;
disk_mem[15737] = 0;
disk_mem[15738] = 0;
disk_mem[15739] = 0;
disk_mem[15740] = 0;
disk_mem[15741] = 0;
disk_mem[15742] = 0;
disk_mem[15743] = 0;
disk_mem[15744] = 0;
disk_mem[15745] = 0;
disk_mem[15746] = 0;
disk_mem[15747] = 0;
disk_mem[15748] = 0;
disk_mem[15749] = 0;
disk_mem[15750] = 0;
disk_mem[15751] = 0;
disk_mem[15752] = 0;
disk_mem[15753] = 0;
disk_mem[15754] = 0;
disk_mem[15755] = 0;
disk_mem[15756] = 0;
disk_mem[15757] = 0;
disk_mem[15758] = 0;
disk_mem[15759] = 0;
disk_mem[15760] = 0;
disk_mem[15761] = 0;
disk_mem[15762] = 0;
disk_mem[15763] = 0;
disk_mem[15764] = 0;
disk_mem[15765] = 0;
disk_mem[15766] = 0;
disk_mem[15767] = 0;
disk_mem[15768] = 0;
disk_mem[15769] = 0;
disk_mem[15770] = 0;
disk_mem[15771] = 0;
disk_mem[15772] = 0;
disk_mem[15773] = 0;
disk_mem[15774] = 0;
disk_mem[15775] = 0;
disk_mem[15776] = 0;
disk_mem[15777] = 0;
disk_mem[15778] = 0;
disk_mem[15779] = 0;
disk_mem[15780] = 0;
disk_mem[15781] = 0;
disk_mem[15782] = 0;
disk_mem[15783] = 0;
disk_mem[15784] = 0;
disk_mem[15785] = 0;
disk_mem[15786] = 0;
disk_mem[15787] = 0;
disk_mem[15788] = 0;
disk_mem[15789] = 0;
disk_mem[15790] = 0;
disk_mem[15791] = 0;
disk_mem[15792] = 0;
disk_mem[15793] = 0;
disk_mem[15794] = 0;
disk_mem[15795] = 0;
disk_mem[15796] = 0;
disk_mem[15797] = 0;
disk_mem[15798] = 0;
disk_mem[15799] = 0;
disk_mem[15800] = 0;
disk_mem[15801] = 0;
disk_mem[15802] = 0;
disk_mem[15803] = 0;
disk_mem[15804] = 0;
disk_mem[15805] = 0;
disk_mem[15806] = 0;
disk_mem[15807] = 0;
disk_mem[15808] = 0;
disk_mem[15809] = 0;
disk_mem[15810] = 0;
disk_mem[15811] = 0;
disk_mem[15812] = 0;
disk_mem[15813] = 0;
disk_mem[15814] = 0;
disk_mem[15815] = 0;
disk_mem[15816] = 0;
disk_mem[15817] = 0;
disk_mem[15818] = 0;
disk_mem[15819] = 0;
disk_mem[15820] = 0;
disk_mem[15821] = 0;
disk_mem[15822] = 0;
disk_mem[15823] = 0;
disk_mem[15824] = 0;
disk_mem[15825] = 0;
disk_mem[15826] = 0;
disk_mem[15827] = 0;
disk_mem[15828] = 0;
disk_mem[15829] = 0;
disk_mem[15830] = 0;
disk_mem[15831] = 0;
disk_mem[15832] = 0;
disk_mem[15833] = 0;
disk_mem[15834] = 0;
disk_mem[15835] = 0;
disk_mem[15836] = 0;
disk_mem[15837] = 0;
disk_mem[15838] = 0;
disk_mem[15839] = 0;
disk_mem[15840] = 0;
disk_mem[15841] = 0;
disk_mem[15842] = 0;
disk_mem[15843] = 0;
disk_mem[15844] = 0;
disk_mem[15845] = 0;
disk_mem[15846] = 0;
disk_mem[15847] = 0;
disk_mem[15848] = 0;
disk_mem[15849] = 0;
disk_mem[15850] = 0;
disk_mem[15851] = 0;
disk_mem[15852] = 0;
disk_mem[15853] = 0;
disk_mem[15854] = 0;
disk_mem[15855] = 0;
disk_mem[15856] = 0;
disk_mem[15857] = 0;
disk_mem[15858] = 0;
disk_mem[15859] = 0;
disk_mem[15860] = 0;
disk_mem[15861] = 0;
disk_mem[15862] = 0;
disk_mem[15863] = 0;
disk_mem[15864] = 0;
disk_mem[15865] = 0;
disk_mem[15866] = 0;
disk_mem[15867] = 0;
disk_mem[15868] = 0;
disk_mem[15869] = 0;
disk_mem[15870] = 0;
disk_mem[15871] = 0;
disk_mem[15872] = 0;
disk_mem[15873] = 0;
disk_mem[15874] = 0;
disk_mem[15875] = 0;
disk_mem[15876] = 0;
disk_mem[15877] = 0;
disk_mem[15878] = 0;
disk_mem[15879] = 0;
disk_mem[15880] = 0;
disk_mem[15881] = 0;
disk_mem[15882] = 0;
disk_mem[15883] = 0;
disk_mem[15884] = 0;
disk_mem[15885] = 0;
disk_mem[15886] = 0;
disk_mem[15887] = 0;
disk_mem[15888] = 0;
disk_mem[15889] = 0;
disk_mem[15890] = 0;
disk_mem[15891] = 0;
disk_mem[15892] = 0;
disk_mem[15893] = 0;
disk_mem[15894] = 0;
disk_mem[15895] = 0;
disk_mem[15896] = 0;
disk_mem[15897] = 0;
disk_mem[15898] = 0;
disk_mem[15899] = 0;
disk_mem[15900] = 0;
disk_mem[15901] = 0;
disk_mem[15902] = 0;
disk_mem[15903] = 0;
disk_mem[15904] = 0;
disk_mem[15905] = 0;
disk_mem[15906] = 0;
disk_mem[15907] = 0;
disk_mem[15908] = 0;
disk_mem[15909] = 0;
disk_mem[15910] = 0;
disk_mem[15911] = 0;
disk_mem[15912] = 0;
disk_mem[15913] = 0;
disk_mem[15914] = 0;
disk_mem[15915] = 0;
disk_mem[15916] = 0;
disk_mem[15917] = 0;
disk_mem[15918] = 0;
disk_mem[15919] = 0;
disk_mem[15920] = 0;
disk_mem[15921] = 0;
disk_mem[15922] = 0;
disk_mem[15923] = 0;
disk_mem[15924] = 0;
disk_mem[15925] = 0;
disk_mem[15926] = 0;
disk_mem[15927] = 0;
disk_mem[15928] = 0;
disk_mem[15929] = 0;
disk_mem[15930] = 0;
disk_mem[15931] = 0;
disk_mem[15932] = 0;
disk_mem[15933] = 0;
disk_mem[15934] = 0;
disk_mem[15935] = 0;
disk_mem[15936] = 0;
disk_mem[15937] = 0;
disk_mem[15938] = 0;
disk_mem[15939] = 0;
disk_mem[15940] = 0;
disk_mem[15941] = 0;
disk_mem[15942] = 0;
disk_mem[15943] = 0;
disk_mem[15944] = 0;
disk_mem[15945] = 0;
disk_mem[15946] = 0;
disk_mem[15947] = 0;
disk_mem[15948] = 0;
disk_mem[15949] = 0;
disk_mem[15950] = 0;
disk_mem[15951] = 0;
disk_mem[15952] = 0;
disk_mem[15953] = 0;
disk_mem[15954] = 0;
disk_mem[15955] = 0;
disk_mem[15956] = 0;
disk_mem[15957] = 0;
disk_mem[15958] = 0;
disk_mem[15959] = 0;
disk_mem[15960] = 0;
disk_mem[15961] = 0;
disk_mem[15962] = 0;
disk_mem[15963] = 0;
disk_mem[15964] = 0;
disk_mem[15965] = 0;
disk_mem[15966] = 0;
disk_mem[15967] = 0;
disk_mem[15968] = 0;
disk_mem[15969] = 0;
disk_mem[15970] = 0;
disk_mem[15971] = 0;
disk_mem[15972] = 0;
disk_mem[15973] = 0;
disk_mem[15974] = 0;
disk_mem[15975] = 0;
disk_mem[15976] = 0;
disk_mem[15977] = 0;
disk_mem[15978] = 0;
disk_mem[15979] = 0;
disk_mem[15980] = 0;
disk_mem[15981] = 0;
disk_mem[15982] = 0;
disk_mem[15983] = 0;
disk_mem[15984] = 0;
disk_mem[15985] = 0;
disk_mem[15986] = 0;
disk_mem[15987] = 0;
disk_mem[15988] = 0;
disk_mem[15989] = 0;
disk_mem[15990] = 0;
disk_mem[15991] = 0;
disk_mem[15992] = 0;
disk_mem[15993] = 0;
disk_mem[15994] = 0;
disk_mem[15995] = 0;
disk_mem[15996] = 0;
disk_mem[15997] = 0;
disk_mem[15998] = 0;
disk_mem[15999] = 0;
disk_mem[16000] = 0;
disk_mem[16001] = 0;
disk_mem[16002] = 0;
disk_mem[16003] = 0;
disk_mem[16004] = 0;
disk_mem[16005] = 0;
disk_mem[16006] = 0;
disk_mem[16007] = 0;
disk_mem[16008] = 0;
disk_mem[16009] = 0;
disk_mem[16010] = 0;
disk_mem[16011] = 0;
disk_mem[16012] = 0;
disk_mem[16013] = 0;
disk_mem[16014] = 0;
disk_mem[16015] = 0;
disk_mem[16016] = 0;
disk_mem[16017] = 0;
disk_mem[16018] = 0;
disk_mem[16019] = 0;
disk_mem[16020] = 0;
disk_mem[16021] = 0;
disk_mem[16022] = 0;
disk_mem[16023] = 0;
disk_mem[16024] = 0;
disk_mem[16025] = 0;
disk_mem[16026] = 0;
disk_mem[16027] = 0;
disk_mem[16028] = 0;
disk_mem[16029] = 0;
disk_mem[16030] = 0;
disk_mem[16031] = 0;
disk_mem[16032] = 0;
disk_mem[16033] = 0;
disk_mem[16034] = 0;
disk_mem[16035] = 0;
disk_mem[16036] = 0;
disk_mem[16037] = 0;
disk_mem[16038] = 0;
disk_mem[16039] = 0;
disk_mem[16040] = 0;
disk_mem[16041] = 0;
disk_mem[16042] = 0;
disk_mem[16043] = 0;
disk_mem[16044] = 0;
disk_mem[16045] = 0;
disk_mem[16046] = 0;
disk_mem[16047] = 0;
disk_mem[16048] = 0;
disk_mem[16049] = 0;
disk_mem[16050] = 0;
disk_mem[16051] = 0;
disk_mem[16052] = 0;
disk_mem[16053] = 0;
disk_mem[16054] = 0;
disk_mem[16055] = 0;
disk_mem[16056] = 0;
disk_mem[16057] = 0;
disk_mem[16058] = 0;
disk_mem[16059] = 0;
disk_mem[16060] = 0;
disk_mem[16061] = 0;
disk_mem[16062] = 0;
disk_mem[16063] = 0;
disk_mem[16064] = 0;
disk_mem[16065] = 0;
disk_mem[16066] = 0;
disk_mem[16067] = 0;
disk_mem[16068] = 0;
disk_mem[16069] = 0;
disk_mem[16070] = 0;
disk_mem[16071] = 0;
disk_mem[16072] = 0;
disk_mem[16073] = 0;
disk_mem[16074] = 0;
disk_mem[16075] = 0;
disk_mem[16076] = 0;
disk_mem[16077] = 0;
disk_mem[16078] = 0;
disk_mem[16079] = 0;
disk_mem[16080] = 0;
disk_mem[16081] = 0;
disk_mem[16082] = 0;
disk_mem[16083] = 0;
disk_mem[16084] = 0;
disk_mem[16085] = 0;
disk_mem[16086] = 0;
disk_mem[16087] = 0;
disk_mem[16088] = 0;
disk_mem[16089] = 0;
disk_mem[16090] = 0;
disk_mem[16091] = 0;
disk_mem[16092] = 0;
disk_mem[16093] = 0;
disk_mem[16094] = 0;
disk_mem[16095] = 0;
disk_mem[16096] = 0;
disk_mem[16097] = 0;
disk_mem[16098] = 0;
disk_mem[16099] = 0;
disk_mem[16100] = 0;
disk_mem[16101] = 0;
disk_mem[16102] = 0;
disk_mem[16103] = 0;
disk_mem[16104] = 0;
disk_mem[16105] = 0;
disk_mem[16106] = 0;
disk_mem[16107] = 0;
disk_mem[16108] = 0;
disk_mem[16109] = 0;
disk_mem[16110] = 0;
disk_mem[16111] = 0;
disk_mem[16112] = 0;
disk_mem[16113] = 0;
disk_mem[16114] = 0;
disk_mem[16115] = 0;
disk_mem[16116] = 0;
disk_mem[16117] = 0;
disk_mem[16118] = 0;
disk_mem[16119] = 0;
disk_mem[16120] = 0;
disk_mem[16121] = 0;
disk_mem[16122] = 0;
disk_mem[16123] = 0;
disk_mem[16124] = 0;
disk_mem[16125] = 0;
disk_mem[16126] = 0;
disk_mem[16127] = 0;
disk_mem[16128] = 0;
disk_mem[16129] = 0;
disk_mem[16130] = 0;
disk_mem[16131] = 0;
disk_mem[16132] = 0;
disk_mem[16133] = 0;
disk_mem[16134] = 0;
disk_mem[16135] = 0;
disk_mem[16136] = 0;
disk_mem[16137] = 0;
disk_mem[16138] = 0;
disk_mem[16139] = 0;
disk_mem[16140] = 0;
disk_mem[16141] = 0;
disk_mem[16142] = 0;
disk_mem[16143] = 0;
disk_mem[16144] = 0;
disk_mem[16145] = 0;
disk_mem[16146] = 0;
disk_mem[16147] = 0;
disk_mem[16148] = 0;
disk_mem[16149] = 0;
disk_mem[16150] = 0;
disk_mem[16151] = 0;
disk_mem[16152] = 0;
disk_mem[16153] = 0;
disk_mem[16154] = 0;
disk_mem[16155] = 0;
disk_mem[16156] = 0;
disk_mem[16157] = 0;
disk_mem[16158] = 0;
disk_mem[16159] = 0;
disk_mem[16160] = 0;
disk_mem[16161] = 0;
disk_mem[16162] = 0;
disk_mem[16163] = 0;
disk_mem[16164] = 0;
disk_mem[16165] = 0;
disk_mem[16166] = 0;
disk_mem[16167] = 0;
disk_mem[16168] = 0;
disk_mem[16169] = 0;
disk_mem[16170] = 0;
disk_mem[16171] = 0;
disk_mem[16172] = 0;
disk_mem[16173] = 0;
disk_mem[16174] = 0;
disk_mem[16175] = 0;
disk_mem[16176] = 0;
disk_mem[16177] = 0;
disk_mem[16178] = 0;
disk_mem[16179] = 0;
disk_mem[16180] = 0;
disk_mem[16181] = 0;
disk_mem[16182] = 0;
disk_mem[16183] = 0;
disk_mem[16184] = 0;
disk_mem[16185] = 0;
disk_mem[16186] = 0;
disk_mem[16187] = 0;
disk_mem[16188] = 0;
disk_mem[16189] = 0;
disk_mem[16190] = 0;
disk_mem[16191] = 0;
disk_mem[16192] = 0;
disk_mem[16193] = 0;
disk_mem[16194] = 0;
disk_mem[16195] = 0;
disk_mem[16196] = 0;
disk_mem[16197] = 0;
disk_mem[16198] = 0;
disk_mem[16199] = 0;
disk_mem[16200] = 0;
disk_mem[16201] = 0;
disk_mem[16202] = 0;
disk_mem[16203] = 0;
disk_mem[16204] = 0;
disk_mem[16205] = 0;
disk_mem[16206] = 0;
disk_mem[16207] = 0;
disk_mem[16208] = 0;
disk_mem[16209] = 0;
disk_mem[16210] = 0;
disk_mem[16211] = 0;
disk_mem[16212] = 0;
disk_mem[16213] = 0;
disk_mem[16214] = 0;
disk_mem[16215] = 0;
disk_mem[16216] = 0;
disk_mem[16217] = 0;
disk_mem[16218] = 0;
disk_mem[16219] = 0;
disk_mem[16220] = 0;
disk_mem[16221] = 0;
disk_mem[16222] = 0;
disk_mem[16223] = 0;
disk_mem[16224] = 0;
disk_mem[16225] = 0;
disk_mem[16226] = 0;
disk_mem[16227] = 0;
disk_mem[16228] = 0;
disk_mem[16229] = 0;
disk_mem[16230] = 0;
disk_mem[16231] = 0;
disk_mem[16232] = 0;
disk_mem[16233] = 0;
disk_mem[16234] = 0;
disk_mem[16235] = 0;
disk_mem[16236] = 0;
disk_mem[16237] = 0;
disk_mem[16238] = 0;
disk_mem[16239] = 0;
disk_mem[16240] = 0;
disk_mem[16241] = 0;
disk_mem[16242] = 0;
disk_mem[16243] = 0;
disk_mem[16244] = 0;
disk_mem[16245] = 0;
disk_mem[16246] = 0;
disk_mem[16247] = 0;
disk_mem[16248] = 0;
disk_mem[16249] = 0;
disk_mem[16250] = 0;
disk_mem[16251] = 0;
disk_mem[16252] = 0;
disk_mem[16253] = 0;
disk_mem[16254] = 0;
disk_mem[16255] = 0;
disk_mem[16256] = 0;
disk_mem[16257] = 0;
disk_mem[16258] = 0;
disk_mem[16259] = 0;
disk_mem[16260] = 0;
disk_mem[16261] = 0;
disk_mem[16262] = 0;
disk_mem[16263] = 0;
disk_mem[16264] = 0;
disk_mem[16265] = 0;
disk_mem[16266] = 0;
disk_mem[16267] = 0;
disk_mem[16268] = 0;
disk_mem[16269] = 0;
disk_mem[16270] = 0;
disk_mem[16271] = 0;
disk_mem[16272] = 0;
disk_mem[16273] = 0;
disk_mem[16274] = 0;
disk_mem[16275] = 0;
disk_mem[16276] = 0;
disk_mem[16277] = 0;
disk_mem[16278] = 0;
disk_mem[16279] = 0;
disk_mem[16280] = 0;
disk_mem[16281] = 0;
disk_mem[16282] = 0;
disk_mem[16283] = 0;
disk_mem[16284] = 0;
disk_mem[16285] = 0;
disk_mem[16286] = 0;
disk_mem[16287] = 0;
disk_mem[16288] = 0;
disk_mem[16289] = 0;
disk_mem[16290] = 0;
disk_mem[16291] = 0;
disk_mem[16292] = 0;
disk_mem[16293] = 0;
disk_mem[16294] = 0;
disk_mem[16295] = 0;
disk_mem[16296] = 0;
disk_mem[16297] = 0;
disk_mem[16298] = 0;
disk_mem[16299] = 0;
disk_mem[16300] = 0;
disk_mem[16301] = 0;
disk_mem[16302] = 0;
disk_mem[16303] = 0;
disk_mem[16304] = 0;
disk_mem[16305] = 0;
disk_mem[16306] = 0;
disk_mem[16307] = 0;
disk_mem[16308] = 0;
disk_mem[16309] = 0;
disk_mem[16310] = 0;
disk_mem[16311] = 0;
disk_mem[16312] = 0;
disk_mem[16313] = 0;
disk_mem[16314] = 0;
disk_mem[16315] = 0;
disk_mem[16316] = 0;
disk_mem[16317] = 0;
disk_mem[16318] = 0;
disk_mem[16319] = 0;
disk_mem[16320] = 0;
disk_mem[16321] = 0;
disk_mem[16322] = 0;
disk_mem[16323] = 0;
disk_mem[16324] = 0;
disk_mem[16325] = 0;
disk_mem[16326] = 0;
disk_mem[16327] = 0;
disk_mem[16328] = 0;
disk_mem[16329] = 0;
disk_mem[16330] = 0;
disk_mem[16331] = 0;
disk_mem[16332] = 0;
disk_mem[16333] = 0;
disk_mem[16334] = 0;
disk_mem[16335] = 0;
disk_mem[16336] = 0;
disk_mem[16337] = 0;
disk_mem[16338] = 0;
disk_mem[16339] = 0;
disk_mem[16340] = 0;
disk_mem[16341] = 0;
disk_mem[16342] = 0;
disk_mem[16343] = 0;
disk_mem[16344] = 0;
disk_mem[16345] = 0;
disk_mem[16346] = 0;
disk_mem[16347] = 0;
disk_mem[16348] = 0;
disk_mem[16349] = 0;
disk_mem[16350] = 0;
disk_mem[16351] = 0;
disk_mem[16352] = 0;
disk_mem[16353] = 0;
disk_mem[16354] = 0;
disk_mem[16355] = 0;
disk_mem[16356] = 0;
disk_mem[16357] = 0;
disk_mem[16358] = 0;
disk_mem[16359] = 0;
disk_mem[16360] = 0;
disk_mem[16361] = 0;
disk_mem[16362] = 0;
disk_mem[16363] = 0;
disk_mem[16364] = 0;
disk_mem[16365] = 0;
disk_mem[16366] = 0;
disk_mem[16367] = 0;
disk_mem[16368] = 0;
disk_mem[16369] = 0;
disk_mem[16370] = 0;
disk_mem[16371] = 0;
disk_mem[16372] = 0;
disk_mem[16373] = 0;
disk_mem[16374] = 0;
disk_mem[16375] = 0;
disk_mem[16376] = 0;
disk_mem[16377] = 0;
disk_mem[16378] = 0;
disk_mem[16379] = 0;
disk_mem[16380] = 0;
disk_mem[16381] = 0;
disk_mem[16382] = 0;
disk_mem[16383] = 0;
disk_mem[16384] = 0;
disk_mem[16385] = 0;
disk_mem[16386] = 0;
disk_mem[16387] = 0;
disk_mem[16388] = 0;
disk_mem[16389] = 0;
disk_mem[16390] = 0;
disk_mem[16391] = 0;
disk_mem[16392] = 0;
disk_mem[16393] = 0;
disk_mem[16394] = 0;
disk_mem[16395] = 0;
disk_mem[16396] = 0;
disk_mem[16397] = 0;
disk_mem[16398] = 0;
disk_mem[16399] = 0;
disk_mem[16400] = 0;
disk_mem[16401] = 0;
disk_mem[16402] = 0;
disk_mem[16403] = 0;
disk_mem[16404] = 0;
disk_mem[16405] = 0;
disk_mem[16406] = 0;
disk_mem[16407] = 0;
disk_mem[16408] = 0;
disk_mem[16409] = 0;
disk_mem[16410] = 0;
disk_mem[16411] = 0;
disk_mem[16412] = 0;
disk_mem[16413] = 0;
disk_mem[16414] = 0;
disk_mem[16415] = 0;
disk_mem[16416] = 0;
disk_mem[16417] = 0;
disk_mem[16418] = 0;
disk_mem[16419] = 0;
disk_mem[16420] = 0;
disk_mem[16421] = 0;
disk_mem[16422] = 0;
disk_mem[16423] = 0;
disk_mem[16424] = 0;
disk_mem[16425] = 0;
disk_mem[16426] = 0;
disk_mem[16427] = 0;
disk_mem[16428] = 0;
disk_mem[16429] = 0;
disk_mem[16430] = 0;
disk_mem[16431] = 0;
disk_mem[16432] = 0;
disk_mem[16433] = 0;
disk_mem[16434] = 0;
disk_mem[16435] = 0;
disk_mem[16436] = 0;
disk_mem[16437] = 0;
disk_mem[16438] = 0;
disk_mem[16439] = 0;
disk_mem[16440] = 0;
disk_mem[16441] = 0;
disk_mem[16442] = 0;
disk_mem[16443] = 0;
disk_mem[16444] = 0;
disk_mem[16445] = 0;
disk_mem[16446] = 0;
disk_mem[16447] = 0;
disk_mem[16448] = 0;
disk_mem[16449] = 0;
disk_mem[16450] = 0;
disk_mem[16451] = 0;
disk_mem[16452] = 0;
disk_mem[16453] = 0;
disk_mem[16454] = 0;
disk_mem[16455] = 0;
disk_mem[16456] = 0;
disk_mem[16457] = 0;
disk_mem[16458] = 0;
disk_mem[16459] = 0;
disk_mem[16460] = 0;
disk_mem[16461] = 0;
disk_mem[16462] = 0;
disk_mem[16463] = 0;
disk_mem[16464] = 0;
disk_mem[16465] = 0;
disk_mem[16466] = 0;
disk_mem[16467] = 0;
disk_mem[16468] = 0;
disk_mem[16469] = 0;
disk_mem[16470] = 0;
disk_mem[16471] = 0;
disk_mem[16472] = 0;
disk_mem[16473] = 0;
disk_mem[16474] = 0;
disk_mem[16475] = 0;
disk_mem[16476] = 0;
disk_mem[16477] = 0;
disk_mem[16478] = 0;
disk_mem[16479] = 0;
disk_mem[16480] = 0;
disk_mem[16481] = 0;
disk_mem[16482] = 0;
disk_mem[16483] = 0;
disk_mem[16484] = 0;
disk_mem[16485] = 0;
disk_mem[16486] = 0;
disk_mem[16487] = 0;
disk_mem[16488] = 0;
disk_mem[16489] = 0;
disk_mem[16490] = 0;
disk_mem[16491] = 0;
disk_mem[16492] = 0;
disk_mem[16493] = 0;
disk_mem[16494] = 0;
disk_mem[16495] = 0;
disk_mem[16496] = 0;
disk_mem[16497] = 0;
disk_mem[16498] = 0;
disk_mem[16499] = 0;
disk_mem[16500] = 0;
disk_mem[16501] = 0;
disk_mem[16502] = 0;
disk_mem[16503] = 0;
disk_mem[16504] = 0;
disk_mem[16505] = 0;
disk_mem[16506] = 0;
disk_mem[16507] = 0;
disk_mem[16508] = 0;
disk_mem[16509] = 0;
disk_mem[16510] = 0;
disk_mem[16511] = 0;
disk_mem[16512] = 0;
disk_mem[16513] = 0;
disk_mem[16514] = 0;
disk_mem[16515] = 0;
disk_mem[16516] = 0;
disk_mem[16517] = 0;
disk_mem[16518] = 0;
disk_mem[16519] = 0;
disk_mem[16520] = 0;
disk_mem[16521] = 0;
disk_mem[16522] = 0;
disk_mem[16523] = 0;
disk_mem[16524] = 0;
disk_mem[16525] = 0;
disk_mem[16526] = 0;
disk_mem[16527] = 0;
disk_mem[16528] = 0;
disk_mem[16529] = 0;
disk_mem[16530] = 0;
disk_mem[16531] = 0;
disk_mem[16532] = 0;
disk_mem[16533] = 0;
disk_mem[16534] = 0;
disk_mem[16535] = 0;
disk_mem[16536] = 0;
disk_mem[16537] = 0;
disk_mem[16538] = 0;
disk_mem[16539] = 0;
disk_mem[16540] = 0;
disk_mem[16541] = 0;
disk_mem[16542] = 0;
disk_mem[16543] = 0;
disk_mem[16544] = 0;
disk_mem[16545] = 0;
disk_mem[16546] = 0;
disk_mem[16547] = 0;
disk_mem[16548] = 0;
disk_mem[16549] = 0;
disk_mem[16550] = 0;
disk_mem[16551] = 0;
disk_mem[16552] = 0;
disk_mem[16553] = 0;
disk_mem[16554] = 0;
disk_mem[16555] = 0;
disk_mem[16556] = 0;
disk_mem[16557] = 0;
disk_mem[16558] = 0;
disk_mem[16559] = 0;
disk_mem[16560] = 0;
disk_mem[16561] = 0;
disk_mem[16562] = 0;
disk_mem[16563] = 0;
disk_mem[16564] = 0;
disk_mem[16565] = 0;
disk_mem[16566] = 0;
disk_mem[16567] = 0;
disk_mem[16568] = 0;
disk_mem[16569] = 0;
disk_mem[16570] = 0;
disk_mem[16571] = 0;
disk_mem[16572] = 0;
disk_mem[16573] = 0;
disk_mem[16574] = 0;
disk_mem[16575] = 0;
disk_mem[16576] = 0;
disk_mem[16577] = 0;
disk_mem[16578] = 0;
disk_mem[16579] = 0;
disk_mem[16580] = 0;
disk_mem[16581] = 0;
disk_mem[16582] = 0;
disk_mem[16583] = 0;
disk_mem[16584] = 0;
disk_mem[16585] = 0;
disk_mem[16586] = 0;
disk_mem[16587] = 0;
disk_mem[16588] = 0;
disk_mem[16589] = 0;
disk_mem[16590] = 0;
disk_mem[16591] = 0;
disk_mem[16592] = 0;
disk_mem[16593] = 0;
disk_mem[16594] = 0;
disk_mem[16595] = 0;
disk_mem[16596] = 0;
disk_mem[16597] = 0;
disk_mem[16598] = 0;
disk_mem[16599] = 0;
disk_mem[16600] = 0;
disk_mem[16601] = 0;
disk_mem[16602] = 0;
disk_mem[16603] = 0;
disk_mem[16604] = 0;
disk_mem[16605] = 0;
disk_mem[16606] = 0;
disk_mem[16607] = 0;
disk_mem[16608] = 0;
disk_mem[16609] = 0;
disk_mem[16610] = 0;
disk_mem[16611] = 0;
disk_mem[16612] = 0;
disk_mem[16613] = 0;
disk_mem[16614] = 0;
disk_mem[16615] = 0;
disk_mem[16616] = 0;
disk_mem[16617] = 0;
disk_mem[16618] = 0;
disk_mem[16619] = 0;
disk_mem[16620] = 0;
disk_mem[16621] = 0;
disk_mem[16622] = 0;
disk_mem[16623] = 0;
disk_mem[16624] = 0;
disk_mem[16625] = 0;
disk_mem[16626] = 0;
disk_mem[16627] = 0;
disk_mem[16628] = 0;
disk_mem[16629] = 0;
disk_mem[16630] = 0;
disk_mem[16631] = 0;
disk_mem[16632] = 0;
disk_mem[16633] = 0;
disk_mem[16634] = 0;
disk_mem[16635] = 0;
disk_mem[16636] = 0;
disk_mem[16637] = 0;
disk_mem[16638] = 0;
disk_mem[16639] = 0;
disk_mem[16640] = 0;
disk_mem[16641] = 0;
disk_mem[16642] = 0;
disk_mem[16643] = 0;
disk_mem[16644] = 0;
disk_mem[16645] = 0;
disk_mem[16646] = 0;
disk_mem[16647] = 0;
disk_mem[16648] = 0;
disk_mem[16649] = 0;
disk_mem[16650] = 0;
disk_mem[16651] = 0;
disk_mem[16652] = 0;
disk_mem[16653] = 0;
disk_mem[16654] = 0;
disk_mem[16655] = 0;
disk_mem[16656] = 0;
disk_mem[16657] = 0;
disk_mem[16658] = 0;
disk_mem[16659] = 0;
disk_mem[16660] = 0;
disk_mem[16661] = 0;
disk_mem[16662] = 0;
disk_mem[16663] = 0;
disk_mem[16664] = 0;
disk_mem[16665] = 0;
disk_mem[16666] = 0;
disk_mem[16667] = 0;
disk_mem[16668] = 0;
disk_mem[16669] = 0;
disk_mem[16670] = 0;
disk_mem[16671] = 0;
disk_mem[16672] = 0;
disk_mem[16673] = 0;
disk_mem[16674] = 0;
disk_mem[16675] = 0;
disk_mem[16676] = 0;
disk_mem[16677] = 0;
disk_mem[16678] = 0;
disk_mem[16679] = 0;
disk_mem[16680] = 0;
disk_mem[16681] = 0;
disk_mem[16682] = 0;
disk_mem[16683] = 0;
disk_mem[16684] = 0;
disk_mem[16685] = 0;
disk_mem[16686] = 0;
disk_mem[16687] = 0;
disk_mem[16688] = 0;
disk_mem[16689] = 0;
disk_mem[16690] = 0;
disk_mem[16691] = 0;
disk_mem[16692] = 0;
disk_mem[16693] = 0;
disk_mem[16694] = 0;
disk_mem[16695] = 0;
disk_mem[16696] = 0;
disk_mem[16697] = 0;
disk_mem[16698] = 0;
disk_mem[16699] = 0;
disk_mem[16700] = 0;
disk_mem[16701] = 0;
disk_mem[16702] = 0;
disk_mem[16703] = 0;
disk_mem[16704] = 0;
disk_mem[16705] = 0;
disk_mem[16706] = 0;
disk_mem[16707] = 0;
disk_mem[16708] = 0;
disk_mem[16709] = 0;
disk_mem[16710] = 0;
disk_mem[16711] = 0;
disk_mem[16712] = 0;
disk_mem[16713] = 0;
disk_mem[16714] = 0;
disk_mem[16715] = 0;
disk_mem[16716] = 0;
disk_mem[16717] = 0;
disk_mem[16718] = 0;
disk_mem[16719] = 0;
disk_mem[16720] = 0;
disk_mem[16721] = 0;
disk_mem[16722] = 0;
disk_mem[16723] = 0;
disk_mem[16724] = 0;
disk_mem[16725] = 0;
disk_mem[16726] = 0;
disk_mem[16727] = 0;
disk_mem[16728] = 0;
disk_mem[16729] = 0;
disk_mem[16730] = 0;
disk_mem[16731] = 0;
disk_mem[16732] = 0;
disk_mem[16733] = 0;
disk_mem[16734] = 0;
disk_mem[16735] = 0;
disk_mem[16736] = 0;
disk_mem[16737] = 0;
disk_mem[16738] = 0;
disk_mem[16739] = 0;
disk_mem[16740] = 0;
disk_mem[16741] = 0;
disk_mem[16742] = 0;
disk_mem[16743] = 0;
disk_mem[16744] = 0;
disk_mem[16745] = 0;
disk_mem[16746] = 0;
disk_mem[16747] = 0;
disk_mem[16748] = 0;
disk_mem[16749] = 0;
disk_mem[16750] = 0;
disk_mem[16751] = 0;
disk_mem[16752] = 0;
disk_mem[16753] = 0;
disk_mem[16754] = 0;
disk_mem[16755] = 0;
disk_mem[16756] = 0;
disk_mem[16757] = 0;
disk_mem[16758] = 0;
disk_mem[16759] = 0;
disk_mem[16760] = 0;
disk_mem[16761] = 0;
disk_mem[16762] = 0;
disk_mem[16763] = 0;
disk_mem[16764] = 0;
disk_mem[16765] = 0;
disk_mem[16766] = 0;
disk_mem[16767] = 0;
disk_mem[16768] = 0;
disk_mem[16769] = 0;
disk_mem[16770] = 0;
disk_mem[16771] = 0;
disk_mem[16772] = 0;
disk_mem[16773] = 0;
disk_mem[16774] = 0;
disk_mem[16775] = 0;
disk_mem[16776] = 0;
disk_mem[16777] = 0;
disk_mem[16778] = 0;
disk_mem[16779] = 0;
disk_mem[16780] = 0;
disk_mem[16781] = 0;
disk_mem[16782] = 0;
disk_mem[16783] = 0;
disk_mem[16784] = 0;
disk_mem[16785] = 0;
disk_mem[16786] = 0;
disk_mem[16787] = 0;
disk_mem[16788] = 0;
disk_mem[16789] = 0;
disk_mem[16790] = 0;
disk_mem[16791] = 0;
disk_mem[16792] = 0;
disk_mem[16793] = 0;
disk_mem[16794] = 0;
disk_mem[16795] = 0;
disk_mem[16796] = 0;
disk_mem[16797] = 0;
disk_mem[16798] = 0;
disk_mem[16799] = 0;
disk_mem[16800] = 0;
disk_mem[16801] = 0;
disk_mem[16802] = 0;
disk_mem[16803] = 0;
disk_mem[16804] = 0;
disk_mem[16805] = 0;
disk_mem[16806] = 0;
disk_mem[16807] = 0;
disk_mem[16808] = 0;
disk_mem[16809] = 0;
disk_mem[16810] = 0;
disk_mem[16811] = 0;
disk_mem[16812] = 0;
disk_mem[16813] = 0;
disk_mem[16814] = 0;
disk_mem[16815] = 0;
disk_mem[16816] = 0;
disk_mem[16817] = 0;
disk_mem[16818] = 0;
disk_mem[16819] = 0;
disk_mem[16820] = 0;
disk_mem[16821] = 0;
disk_mem[16822] = 0;
disk_mem[16823] = 0;
disk_mem[16824] = 0;
disk_mem[16825] = 0;
disk_mem[16826] = 0;
disk_mem[16827] = 0;
disk_mem[16828] = 0;
disk_mem[16829] = 0;
disk_mem[16830] = 0;
disk_mem[16831] = 0;
disk_mem[16832] = 0;
disk_mem[16833] = 0;
disk_mem[16834] = 0;
disk_mem[16835] = 0;
disk_mem[16836] = 0;
disk_mem[16837] = 0;
disk_mem[16838] = 0;
disk_mem[16839] = 0;
disk_mem[16840] = 0;
disk_mem[16841] = 0;
disk_mem[16842] = 0;
disk_mem[16843] = 0;
disk_mem[16844] = 0;
disk_mem[16845] = 0;
disk_mem[16846] = 0;
disk_mem[16847] = 0;
disk_mem[16848] = 0;
disk_mem[16849] = 0;
disk_mem[16850] = 0;
disk_mem[16851] = 0;
disk_mem[16852] = 0;
disk_mem[16853] = 0;
disk_mem[16854] = 0;
disk_mem[16855] = 0;
disk_mem[16856] = 0;
disk_mem[16857] = 0;
disk_mem[16858] = 0;
disk_mem[16859] = 0;
disk_mem[16860] = 0;
disk_mem[16861] = 0;
disk_mem[16862] = 0;
disk_mem[16863] = 0;
disk_mem[16864] = 0;
disk_mem[16865] = 0;
disk_mem[16866] = 0;
disk_mem[16867] = 0;
disk_mem[16868] = 0;
disk_mem[16869] = 0;
disk_mem[16870] = 0;
disk_mem[16871] = 0;
disk_mem[16872] = 0;
disk_mem[16873] = 0;
disk_mem[16874] = 0;
disk_mem[16875] = 0;
disk_mem[16876] = 0;
disk_mem[16877] = 0;
disk_mem[16878] = 0;
disk_mem[16879] = 0;
disk_mem[16880] = 0;
disk_mem[16881] = 0;
disk_mem[16882] = 0;
disk_mem[16883] = 0;
disk_mem[16884] = 0;
disk_mem[16885] = 0;
disk_mem[16886] = 0;
disk_mem[16887] = 0;
disk_mem[16888] = 0;
disk_mem[16889] = 0;
disk_mem[16890] = 0;
disk_mem[16891] = 0;
disk_mem[16892] = 0;
disk_mem[16893] = 0;
disk_mem[16894] = 0;
disk_mem[16895] = 0;
disk_mem[16896] = 0;
disk_mem[16897] = 0;
disk_mem[16898] = 0;
disk_mem[16899] = 0;
disk_mem[16900] = 0;
disk_mem[16901] = 0;
disk_mem[16902] = 0;
disk_mem[16903] = 0;
disk_mem[16904] = 0;
disk_mem[16905] = 0;
disk_mem[16906] = 0;
disk_mem[16907] = 0;
disk_mem[16908] = 0;
disk_mem[16909] = 0;
disk_mem[16910] = 0;
disk_mem[16911] = 0;
disk_mem[16912] = 0;
disk_mem[16913] = 0;
disk_mem[16914] = 0;
disk_mem[16915] = 0;
disk_mem[16916] = 0;
disk_mem[16917] = 0;
disk_mem[16918] = 0;
disk_mem[16919] = 0;
disk_mem[16920] = 0;
disk_mem[16921] = 0;
disk_mem[16922] = 0;
disk_mem[16923] = 0;
disk_mem[16924] = 0;
disk_mem[16925] = 0;
disk_mem[16926] = 0;
disk_mem[16927] = 0;
disk_mem[16928] = 0;
disk_mem[16929] = 0;
disk_mem[16930] = 0;
disk_mem[16931] = 0;
disk_mem[16932] = 0;
disk_mem[16933] = 0;
disk_mem[16934] = 0;
disk_mem[16935] = 0;
disk_mem[16936] = 0;
disk_mem[16937] = 0;
disk_mem[16938] = 0;
disk_mem[16939] = 0;
disk_mem[16940] = 0;
disk_mem[16941] = 0;
disk_mem[16942] = 0;
disk_mem[16943] = 0;
disk_mem[16944] = 0;
disk_mem[16945] = 0;
disk_mem[16946] = 0;
disk_mem[16947] = 0;
disk_mem[16948] = 0;
disk_mem[16949] = 0;
disk_mem[16950] = 0;
disk_mem[16951] = 0;
disk_mem[16952] = 0;
disk_mem[16953] = 0;
disk_mem[16954] = 0;
disk_mem[16955] = 0;
disk_mem[16956] = 0;
disk_mem[16957] = 0;
disk_mem[16958] = 0;
disk_mem[16959] = 0;
disk_mem[16960] = 0;
disk_mem[16961] = 0;
disk_mem[16962] = 0;
disk_mem[16963] = 0;
disk_mem[16964] = 0;
disk_mem[16965] = 0;
disk_mem[16966] = 0;
disk_mem[16967] = 0;
disk_mem[16968] = 0;
disk_mem[16969] = 0;
disk_mem[16970] = 0;
disk_mem[16971] = 0;
disk_mem[16972] = 0;
disk_mem[16973] = 0;
disk_mem[16974] = 0;
disk_mem[16975] = 0;
disk_mem[16976] = 0;
disk_mem[16977] = 0;
disk_mem[16978] = 0;
disk_mem[16979] = 0;
disk_mem[16980] = 0;
disk_mem[16981] = 0;
disk_mem[16982] = 0;
disk_mem[16983] = 0;
disk_mem[16984] = 0;
disk_mem[16985] = 0;
disk_mem[16986] = 0;
disk_mem[16987] = 0;
disk_mem[16988] = 0;
disk_mem[16989] = 0;
disk_mem[16990] = 0;
disk_mem[16991] = 0;
disk_mem[16992] = 0;
disk_mem[16993] = 0;
disk_mem[16994] = 0;
disk_mem[16995] = 0;
disk_mem[16996] = 0;
disk_mem[16997] = 0;
disk_mem[16998] = 0;
disk_mem[16999] = 0;
disk_mem[17000] = 0;
disk_mem[17001] = 0;
disk_mem[17002] = 0;
disk_mem[17003] = 0;
disk_mem[17004] = 0;
disk_mem[17005] = 0;
disk_mem[17006] = 0;
disk_mem[17007] = 0;
disk_mem[17008] = 0;
disk_mem[17009] = 0;
disk_mem[17010] = 0;
disk_mem[17011] = 0;
disk_mem[17012] = 0;
disk_mem[17013] = 0;
disk_mem[17014] = 0;
disk_mem[17015] = 0;
disk_mem[17016] = 0;
disk_mem[17017] = 0;
disk_mem[17018] = 0;
disk_mem[17019] = 0;
disk_mem[17020] = 0;
disk_mem[17021] = 0;
disk_mem[17022] = 0;
disk_mem[17023] = 0;
disk_mem[17024] = 0;
disk_mem[17025] = 0;
disk_mem[17026] = 0;
disk_mem[17027] = 0;
disk_mem[17028] = 0;
disk_mem[17029] = 0;
disk_mem[17030] = 0;
disk_mem[17031] = 0;
disk_mem[17032] = 0;
disk_mem[17033] = 0;
disk_mem[17034] = 0;
disk_mem[17035] = 0;
disk_mem[17036] = 0;
disk_mem[17037] = 0;
disk_mem[17038] = 0;
disk_mem[17039] = 0;
disk_mem[17040] = 0;
disk_mem[17041] = 0;
disk_mem[17042] = 0;
disk_mem[17043] = 0;
disk_mem[17044] = 0;
disk_mem[17045] = 0;
disk_mem[17046] = 0;
disk_mem[17047] = 0;
disk_mem[17048] = 0;
disk_mem[17049] = 0;
disk_mem[17050] = 0;
disk_mem[17051] = 0;
disk_mem[17052] = 0;
disk_mem[17053] = 0;
disk_mem[17054] = 0;
disk_mem[17055] = 0;
disk_mem[17056] = 0;
disk_mem[17057] = 0;
disk_mem[17058] = 0;
disk_mem[17059] = 0;
disk_mem[17060] = 0;
disk_mem[17061] = 0;
disk_mem[17062] = 0;
disk_mem[17063] = 0;
disk_mem[17064] = 0;
disk_mem[17065] = 0;
disk_mem[17066] = 0;
disk_mem[17067] = 0;
disk_mem[17068] = 0;
disk_mem[17069] = 0;
disk_mem[17070] = 0;
disk_mem[17071] = 0;
disk_mem[17072] = 0;
disk_mem[17073] = 0;
disk_mem[17074] = 0;
disk_mem[17075] = 0;
disk_mem[17076] = 0;
disk_mem[17077] = 0;
disk_mem[17078] = 0;
disk_mem[17079] = 0;
disk_mem[17080] = 0;
disk_mem[17081] = 0;
disk_mem[17082] = 0;
disk_mem[17083] = 0;
disk_mem[17084] = 0;
disk_mem[17085] = 0;
disk_mem[17086] = 0;
disk_mem[17087] = 0;
disk_mem[17088] = 0;
disk_mem[17089] = 0;
disk_mem[17090] = 0;
disk_mem[17091] = 0;
disk_mem[17092] = 0;
disk_mem[17093] = 0;
disk_mem[17094] = 0;
disk_mem[17095] = 0;
disk_mem[17096] = 0;
disk_mem[17097] = 0;
disk_mem[17098] = 0;
disk_mem[17099] = 0;
disk_mem[17100] = 0;
disk_mem[17101] = 0;
disk_mem[17102] = 0;
disk_mem[17103] = 0;
disk_mem[17104] = 0;
disk_mem[17105] = 0;
disk_mem[17106] = 0;
disk_mem[17107] = 0;
disk_mem[17108] = 0;
disk_mem[17109] = 0;
disk_mem[17110] = 0;
disk_mem[17111] = 0;
disk_mem[17112] = 0;
disk_mem[17113] = 0;
disk_mem[17114] = 0;
disk_mem[17115] = 0;
disk_mem[17116] = 0;
disk_mem[17117] = 0;
disk_mem[17118] = 0;
disk_mem[17119] = 0;
disk_mem[17120] = 0;
disk_mem[17121] = 0;
disk_mem[17122] = 0;
disk_mem[17123] = 0;
disk_mem[17124] = 0;
disk_mem[17125] = 0;
disk_mem[17126] = 0;
disk_mem[17127] = 0;
disk_mem[17128] = 0;
disk_mem[17129] = 0;
disk_mem[17130] = 0;
disk_mem[17131] = 0;
disk_mem[17132] = 0;
disk_mem[17133] = 0;
disk_mem[17134] = 0;
disk_mem[17135] = 0;
disk_mem[17136] = 0;
disk_mem[17137] = 0;
disk_mem[17138] = 0;
disk_mem[17139] = 0;
disk_mem[17140] = 0;
disk_mem[17141] = 0;
disk_mem[17142] = 0;
disk_mem[17143] = 0;
disk_mem[17144] = 0;
disk_mem[17145] = 0;
disk_mem[17146] = 0;
disk_mem[17147] = 0;
disk_mem[17148] = 0;
disk_mem[17149] = 0;
disk_mem[17150] = 0;
disk_mem[17151] = 0;
disk_mem[17152] = 0;
disk_mem[17153] = 0;
disk_mem[17154] = 0;
disk_mem[17155] = 0;
disk_mem[17156] = 0;
disk_mem[17157] = 0;
disk_mem[17158] = 0;
disk_mem[17159] = 0;
disk_mem[17160] = 0;
disk_mem[17161] = 0;
disk_mem[17162] = 0;
disk_mem[17163] = 0;
disk_mem[17164] = 0;
disk_mem[17165] = 0;
disk_mem[17166] = 0;
disk_mem[17167] = 0;
disk_mem[17168] = 0;
disk_mem[17169] = 0;
disk_mem[17170] = 0;
disk_mem[17171] = 0;
disk_mem[17172] = 0;
disk_mem[17173] = 0;
disk_mem[17174] = 0;
disk_mem[17175] = 0;
disk_mem[17176] = 0;
disk_mem[17177] = 0;
disk_mem[17178] = 0;
disk_mem[17179] = 0;
disk_mem[17180] = 0;
disk_mem[17181] = 0;
disk_mem[17182] = 0;
disk_mem[17183] = 0;
disk_mem[17184] = 0;
disk_mem[17185] = 0;
disk_mem[17186] = 0;
disk_mem[17187] = 0;
disk_mem[17188] = 0;
disk_mem[17189] = 0;
disk_mem[17190] = 0;
disk_mem[17191] = 0;
disk_mem[17192] = 0;
disk_mem[17193] = 0;
disk_mem[17194] = 0;
disk_mem[17195] = 0;
disk_mem[17196] = 0;
disk_mem[17197] = 0;
disk_mem[17198] = 0;
disk_mem[17199] = 0;
disk_mem[17200] = 0;
disk_mem[17201] = 0;
disk_mem[17202] = 0;
disk_mem[17203] = 0;
disk_mem[17204] = 0;
disk_mem[17205] = 0;
disk_mem[17206] = 0;
disk_mem[17207] = 0;
disk_mem[17208] = 0;
disk_mem[17209] = 0;
disk_mem[17210] = 0;
disk_mem[17211] = 0;
disk_mem[17212] = 0;
disk_mem[17213] = 0;
disk_mem[17214] = 0;
disk_mem[17215] = 0;
disk_mem[17216] = 0;
disk_mem[17217] = 0;
disk_mem[17218] = 0;
disk_mem[17219] = 0;
disk_mem[17220] = 0;
disk_mem[17221] = 0;
disk_mem[17222] = 0;
disk_mem[17223] = 0;
disk_mem[17224] = 0;
disk_mem[17225] = 0;
disk_mem[17226] = 0;
disk_mem[17227] = 0;
disk_mem[17228] = 0;
disk_mem[17229] = 0;
disk_mem[17230] = 0;
disk_mem[17231] = 0;
disk_mem[17232] = 0;
disk_mem[17233] = 0;
disk_mem[17234] = 0;
disk_mem[17235] = 0;
disk_mem[17236] = 0;
disk_mem[17237] = 0;
disk_mem[17238] = 0;
disk_mem[17239] = 0;
disk_mem[17240] = 0;
disk_mem[17241] = 0;
disk_mem[17242] = 0;
disk_mem[17243] = 0;
disk_mem[17244] = 0;
disk_mem[17245] = 0;
disk_mem[17246] = 0;
disk_mem[17247] = 0;
disk_mem[17248] = 0;
disk_mem[17249] = 0;
disk_mem[17250] = 0;
disk_mem[17251] = 0;
disk_mem[17252] = 0;
disk_mem[17253] = 0;
disk_mem[17254] = 0;
disk_mem[17255] = 0;
disk_mem[17256] = 0;
disk_mem[17257] = 0;
disk_mem[17258] = 0;
disk_mem[17259] = 0;
disk_mem[17260] = 0;
disk_mem[17261] = 0;
disk_mem[17262] = 0;
disk_mem[17263] = 0;
disk_mem[17264] = 0;
disk_mem[17265] = 0;
disk_mem[17266] = 0;
disk_mem[17267] = 0;
disk_mem[17268] = 0;
disk_mem[17269] = 0;
disk_mem[17270] = 0;
disk_mem[17271] = 0;
disk_mem[17272] = 0;
disk_mem[17273] = 0;
disk_mem[17274] = 0;
disk_mem[17275] = 0;
disk_mem[17276] = 0;
disk_mem[17277] = 0;
disk_mem[17278] = 0;
disk_mem[17279] = 0;
disk_mem[17280] = 0;
disk_mem[17281] = 0;
disk_mem[17282] = 0;
disk_mem[17283] = 0;
disk_mem[17284] = 0;
disk_mem[17285] = 0;
disk_mem[17286] = 0;
disk_mem[17287] = 0;
disk_mem[17288] = 0;
disk_mem[17289] = 0;
disk_mem[17290] = 0;
disk_mem[17291] = 0;
disk_mem[17292] = 0;
disk_mem[17293] = 0;
disk_mem[17294] = 0;
disk_mem[17295] = 0;
disk_mem[17296] = 0;
disk_mem[17297] = 0;
disk_mem[17298] = 0;
disk_mem[17299] = 0;
disk_mem[17300] = 0;
disk_mem[17301] = 0;
disk_mem[17302] = 0;
disk_mem[17303] = 0;
disk_mem[17304] = 0;
disk_mem[17305] = 0;
disk_mem[17306] = 0;
disk_mem[17307] = 0;
disk_mem[17308] = 0;
disk_mem[17309] = 0;
disk_mem[17310] = 0;
disk_mem[17311] = 0;
disk_mem[17312] = 0;
disk_mem[17313] = 0;
disk_mem[17314] = 0;
disk_mem[17315] = 0;
disk_mem[17316] = 0;
disk_mem[17317] = 0;
disk_mem[17318] = 0;
disk_mem[17319] = 0;
disk_mem[17320] = 0;
disk_mem[17321] = 0;
disk_mem[17322] = 0;
disk_mem[17323] = 0;
disk_mem[17324] = 0;
disk_mem[17325] = 0;
disk_mem[17326] = 0;
disk_mem[17327] = 0;
disk_mem[17328] = 0;
disk_mem[17329] = 0;
disk_mem[17330] = 0;
disk_mem[17331] = 0;
disk_mem[17332] = 0;
disk_mem[17333] = 0;
disk_mem[17334] = 0;
disk_mem[17335] = 0;
disk_mem[17336] = 0;
disk_mem[17337] = 0;
disk_mem[17338] = 0;
disk_mem[17339] = 0;
disk_mem[17340] = 0;
disk_mem[17341] = 0;
disk_mem[17342] = 0;
disk_mem[17343] = 0;
disk_mem[17344] = 0;
disk_mem[17345] = 0;
disk_mem[17346] = 0;
disk_mem[17347] = 0;
disk_mem[17348] = 0;
disk_mem[17349] = 0;
disk_mem[17350] = 0;
disk_mem[17351] = 0;
disk_mem[17352] = 0;
disk_mem[17353] = 0;
disk_mem[17354] = 0;
disk_mem[17355] = 0;
disk_mem[17356] = 0;
disk_mem[17357] = 0;
disk_mem[17358] = 0;
disk_mem[17359] = 0;
disk_mem[17360] = 0;
disk_mem[17361] = 0;
disk_mem[17362] = 0;
disk_mem[17363] = 0;
disk_mem[17364] = 0;
disk_mem[17365] = 0;
disk_mem[17366] = 0;
disk_mem[17367] = 0;
disk_mem[17368] = 0;
disk_mem[17369] = 0;
disk_mem[17370] = 0;
disk_mem[17371] = 0;
disk_mem[17372] = 0;
disk_mem[17373] = 0;
disk_mem[17374] = 0;
disk_mem[17375] = 0;
disk_mem[17376] = 0;
disk_mem[17377] = 0;
disk_mem[17378] = 0;
disk_mem[17379] = 0;
disk_mem[17380] = 0;
disk_mem[17381] = 0;
disk_mem[17382] = 0;
disk_mem[17383] = 0;
disk_mem[17384] = 0;
disk_mem[17385] = 0;
disk_mem[17386] = 0;
disk_mem[17387] = 0;
disk_mem[17388] = 0;
disk_mem[17389] = 0;
disk_mem[17390] = 0;
disk_mem[17391] = 0;
disk_mem[17392] = 0;
disk_mem[17393] = 0;
disk_mem[17394] = 0;
disk_mem[17395] = 0;
disk_mem[17396] = 0;
disk_mem[17397] = 0;
disk_mem[17398] = 0;
disk_mem[17399] = 0;
disk_mem[17400] = 0;
disk_mem[17401] = 0;
disk_mem[17402] = 0;
disk_mem[17403] = 0;
disk_mem[17404] = 0;
disk_mem[17405] = 0;
disk_mem[17406] = 0;
disk_mem[17407] = 0;
disk_mem[17408] = 0;
disk_mem[17409] = 0;
disk_mem[17410] = 0;
disk_mem[17411] = 0;
disk_mem[17412] = 0;
disk_mem[17413] = 0;
disk_mem[17414] = 0;
disk_mem[17415] = 0;
disk_mem[17416] = 0;
disk_mem[17417] = 0;
disk_mem[17418] = 0;
disk_mem[17419] = 0;
disk_mem[17420] = 0;
disk_mem[17421] = 0;
disk_mem[17422] = 0;
disk_mem[17423] = 0;
disk_mem[17424] = 0;
disk_mem[17425] = 0;
disk_mem[17426] = 0;
disk_mem[17427] = 0;
disk_mem[17428] = 0;
disk_mem[17429] = 0;
disk_mem[17430] = 0;
disk_mem[17431] = 0;
disk_mem[17432] = 0;
disk_mem[17433] = 0;
disk_mem[17434] = 0;
disk_mem[17435] = 0;
disk_mem[17436] = 0;
disk_mem[17437] = 0;
disk_mem[17438] = 0;
disk_mem[17439] = 0;
disk_mem[17440] = 0;
disk_mem[17441] = 0;
disk_mem[17442] = 0;
disk_mem[17443] = 0;
disk_mem[17444] = 0;
disk_mem[17445] = 0;
disk_mem[17446] = 0;
disk_mem[17447] = 0;
disk_mem[17448] = 0;
disk_mem[17449] = 0;
disk_mem[17450] = 0;
disk_mem[17451] = 0;
disk_mem[17452] = 0;
disk_mem[17453] = 0;
disk_mem[17454] = 0;
disk_mem[17455] = 0;
disk_mem[17456] = 0;
disk_mem[17457] = 0;
disk_mem[17458] = 0;
disk_mem[17459] = 0;
disk_mem[17460] = 0;
disk_mem[17461] = 0;
disk_mem[17462] = 0;
disk_mem[17463] = 0;
disk_mem[17464] = 0;
disk_mem[17465] = 0;
disk_mem[17466] = 0;
disk_mem[17467] = 0;
disk_mem[17468] = 0;
disk_mem[17469] = 0;
disk_mem[17470] = 0;
disk_mem[17471] = 0;
disk_mem[17472] = 0;
disk_mem[17473] = 0;
disk_mem[17474] = 0;
disk_mem[17475] = 0;
disk_mem[17476] = 0;
disk_mem[17477] = 0;
disk_mem[17478] = 0;
disk_mem[17479] = 0;
disk_mem[17480] = 0;
disk_mem[17481] = 0;
disk_mem[17482] = 0;
disk_mem[17483] = 0;
disk_mem[17484] = 0;
disk_mem[17485] = 0;
disk_mem[17486] = 0;
disk_mem[17487] = 0;
disk_mem[17488] = 0;
disk_mem[17489] = 0;
disk_mem[17490] = 0;
disk_mem[17491] = 0;
disk_mem[17492] = 0;
disk_mem[17493] = 0;
disk_mem[17494] = 0;
disk_mem[17495] = 0;
disk_mem[17496] = 0;
disk_mem[17497] = 0;
disk_mem[17498] = 0;
disk_mem[17499] = 0;
disk_mem[17500] = 0;
disk_mem[17501] = 0;
disk_mem[17502] = 0;
disk_mem[17503] = 0;
disk_mem[17504] = 0;
disk_mem[17505] = 0;
disk_mem[17506] = 0;
disk_mem[17507] = 0;
disk_mem[17508] = 0;
disk_mem[17509] = 0;
disk_mem[17510] = 0;
disk_mem[17511] = 0;
disk_mem[17512] = 0;
disk_mem[17513] = 0;
disk_mem[17514] = 0;
disk_mem[17515] = 0;
disk_mem[17516] = 0;
disk_mem[17517] = 0;
disk_mem[17518] = 0;
disk_mem[17519] = 0;
disk_mem[17520] = 0;
disk_mem[17521] = 0;
disk_mem[17522] = 0;
disk_mem[17523] = 0;
disk_mem[17524] = 0;
disk_mem[17525] = 0;
disk_mem[17526] = 0;
disk_mem[17527] = 0;
disk_mem[17528] = 0;
disk_mem[17529] = 0;
disk_mem[17530] = 0;
disk_mem[17531] = 0;
disk_mem[17532] = 0;
disk_mem[17533] = 0;
disk_mem[17534] = 0;
disk_mem[17535] = 0;
disk_mem[17536] = 0;
disk_mem[17537] = 0;
disk_mem[17538] = 0;
disk_mem[17539] = 0;
disk_mem[17540] = 0;
disk_mem[17541] = 0;
disk_mem[17542] = 0;
disk_mem[17543] = 0;
disk_mem[17544] = 0;
disk_mem[17545] = 0;
disk_mem[17546] = 0;
disk_mem[17547] = 0;
disk_mem[17548] = 0;
disk_mem[17549] = 0;
disk_mem[17550] = 0;
disk_mem[17551] = 0;
disk_mem[17552] = 0;
disk_mem[17553] = 0;
disk_mem[17554] = 0;
disk_mem[17555] = 0;
disk_mem[17556] = 0;
disk_mem[17557] = 0;
disk_mem[17558] = 0;
disk_mem[17559] = 0;
disk_mem[17560] = 0;
disk_mem[17561] = 0;
disk_mem[17562] = 0;
disk_mem[17563] = 0;
disk_mem[17564] = 0;
disk_mem[17565] = 0;
disk_mem[17566] = 0;
disk_mem[17567] = 0;
disk_mem[17568] = 0;
disk_mem[17569] = 0;
disk_mem[17570] = 0;
disk_mem[17571] = 0;
disk_mem[17572] = 0;
disk_mem[17573] = 0;
disk_mem[17574] = 0;
disk_mem[17575] = 0;
disk_mem[17576] = 0;
disk_mem[17577] = 0;
disk_mem[17578] = 0;
disk_mem[17579] = 0;
disk_mem[17580] = 0;
disk_mem[17581] = 0;
disk_mem[17582] = 0;
disk_mem[17583] = 0;
disk_mem[17584] = 0;
disk_mem[17585] = 0;
disk_mem[17586] = 0;
disk_mem[17587] = 0;
disk_mem[17588] = 0;
disk_mem[17589] = 0;
disk_mem[17590] = 0;
disk_mem[17591] = 0;
disk_mem[17592] = 0;
disk_mem[17593] = 0;
disk_mem[17594] = 0;
disk_mem[17595] = 0;
disk_mem[17596] = 0;
disk_mem[17597] = 0;
disk_mem[17598] = 0;
disk_mem[17599] = 0;
disk_mem[17600] = 0;
disk_mem[17601] = 0;
disk_mem[17602] = 0;
disk_mem[17603] = 0;
disk_mem[17604] = 0;
disk_mem[17605] = 0;
disk_mem[17606] = 0;
disk_mem[17607] = 0;
disk_mem[17608] = 0;
disk_mem[17609] = 0;
disk_mem[17610] = 0;
disk_mem[17611] = 0;
disk_mem[17612] = 0;
disk_mem[17613] = 0;
disk_mem[17614] = 0;
disk_mem[17615] = 0;
disk_mem[17616] = 0;
disk_mem[17617] = 0;
disk_mem[17618] = 0;
disk_mem[17619] = 0;
disk_mem[17620] = 0;
disk_mem[17621] = 0;
disk_mem[17622] = 0;
disk_mem[17623] = 0;
disk_mem[17624] = 0;
disk_mem[17625] = 0;
disk_mem[17626] = 0;
disk_mem[17627] = 0;
disk_mem[17628] = 0;
disk_mem[17629] = 0;
disk_mem[17630] = 0;
disk_mem[17631] = 0;
disk_mem[17632] = 0;
disk_mem[17633] = 0;
disk_mem[17634] = 0;
disk_mem[17635] = 0;
disk_mem[17636] = 0;
disk_mem[17637] = 0;
disk_mem[17638] = 0;
disk_mem[17639] = 0;
disk_mem[17640] = 0;
disk_mem[17641] = 0;
disk_mem[17642] = 0;
disk_mem[17643] = 0;
disk_mem[17644] = 0;
disk_mem[17645] = 0;
disk_mem[17646] = 0;
disk_mem[17647] = 0;
disk_mem[17648] = 0;
disk_mem[17649] = 0;
disk_mem[17650] = 0;
disk_mem[17651] = 0;
disk_mem[17652] = 0;
disk_mem[17653] = 0;
disk_mem[17654] = 0;
disk_mem[17655] = 0;
disk_mem[17656] = 0;
disk_mem[17657] = 0;
disk_mem[17658] = 0;
disk_mem[17659] = 0;
disk_mem[17660] = 0;
disk_mem[17661] = 0;
disk_mem[17662] = 0;
disk_mem[17663] = 0;
disk_mem[17664] = 0;
disk_mem[17665] = 0;
disk_mem[17666] = 0;
disk_mem[17667] = 0;
disk_mem[17668] = 0;
disk_mem[17669] = 0;
disk_mem[17670] = 0;
disk_mem[17671] = 0;
disk_mem[17672] = 0;
disk_mem[17673] = 0;
disk_mem[17674] = 0;
disk_mem[17675] = 0;
disk_mem[17676] = 0;
disk_mem[17677] = 0;
disk_mem[17678] = 0;
disk_mem[17679] = 0;
disk_mem[17680] = 0;
disk_mem[17681] = 0;
disk_mem[17682] = 0;
disk_mem[17683] = 0;
disk_mem[17684] = 0;
disk_mem[17685] = 0;
disk_mem[17686] = 0;
disk_mem[17687] = 0;
disk_mem[17688] = 0;
disk_mem[17689] = 0;
disk_mem[17690] = 0;
disk_mem[17691] = 0;
disk_mem[17692] = 0;
disk_mem[17693] = 0;
disk_mem[17694] = 0;
disk_mem[17695] = 0;
disk_mem[17696] = 0;
disk_mem[17697] = 0;
disk_mem[17698] = 0;
disk_mem[17699] = 0;
disk_mem[17700] = 0;
disk_mem[17701] = 0;
disk_mem[17702] = 0;
disk_mem[17703] = 0;
disk_mem[17704] = 0;
disk_mem[17705] = 0;
disk_mem[17706] = 0;
disk_mem[17707] = 0;
disk_mem[17708] = 0;
disk_mem[17709] = 0;
disk_mem[17710] = 0;
disk_mem[17711] = 0;
disk_mem[17712] = 0;
disk_mem[17713] = 0;
disk_mem[17714] = 0;
disk_mem[17715] = 0;
disk_mem[17716] = 0;
disk_mem[17717] = 0;
disk_mem[17718] = 0;
disk_mem[17719] = 0;
disk_mem[17720] = 0;
disk_mem[17721] = 0;
disk_mem[17722] = 0;
disk_mem[17723] = 0;
disk_mem[17724] = 0;
disk_mem[17725] = 0;
disk_mem[17726] = 0;
disk_mem[17727] = 0;
disk_mem[17728] = 0;
disk_mem[17729] = 0;
disk_mem[17730] = 0;
disk_mem[17731] = 0;
disk_mem[17732] = 0;
disk_mem[17733] = 0;
disk_mem[17734] = 0;
disk_mem[17735] = 0;
disk_mem[17736] = 0;
disk_mem[17737] = 0;
disk_mem[17738] = 0;
disk_mem[17739] = 0;
disk_mem[17740] = 0;
disk_mem[17741] = 0;
disk_mem[17742] = 0;
disk_mem[17743] = 0;
disk_mem[17744] = 0;
disk_mem[17745] = 0;
disk_mem[17746] = 0;
disk_mem[17747] = 0;
disk_mem[17748] = 0;
disk_mem[17749] = 0;
disk_mem[17750] = 0;
disk_mem[17751] = 0;
disk_mem[17752] = 0;
disk_mem[17753] = 0;
disk_mem[17754] = 0;
disk_mem[17755] = 0;
disk_mem[17756] = 0;
disk_mem[17757] = 0;
disk_mem[17758] = 0;
disk_mem[17759] = 0;
disk_mem[17760] = 0;
disk_mem[17761] = 0;
disk_mem[17762] = 0;
disk_mem[17763] = 0;
disk_mem[17764] = 0;
disk_mem[17765] = 0;
disk_mem[17766] = 0;
disk_mem[17767] = 0;
disk_mem[17768] = 0;
disk_mem[17769] = 0;
disk_mem[17770] = 0;
disk_mem[17771] = 0;
disk_mem[17772] = 0;
disk_mem[17773] = 0;
disk_mem[17774] = 0;
disk_mem[17775] = 0;
disk_mem[17776] = 0;
disk_mem[17777] = 0;
disk_mem[17778] = 0;
disk_mem[17779] = 0;
disk_mem[17780] = 0;
disk_mem[17781] = 0;
disk_mem[17782] = 0;
disk_mem[17783] = 0;
disk_mem[17784] = 0;
disk_mem[17785] = 0;
disk_mem[17786] = 0;
disk_mem[17787] = 0;
disk_mem[17788] = 0;
disk_mem[17789] = 0;
disk_mem[17790] = 0;
disk_mem[17791] = 0;
disk_mem[17792] = 0;
disk_mem[17793] = 0;
disk_mem[17794] = 0;
disk_mem[17795] = 0;
disk_mem[17796] = 0;
disk_mem[17797] = 0;
disk_mem[17798] = 0;
disk_mem[17799] = 0;
disk_mem[17800] = 0;
disk_mem[17801] = 0;
disk_mem[17802] = 0;
disk_mem[17803] = 0;
disk_mem[17804] = 0;
disk_mem[17805] = 0;
disk_mem[17806] = 0;
disk_mem[17807] = 0;
disk_mem[17808] = 0;
disk_mem[17809] = 0;
disk_mem[17810] = 0;
disk_mem[17811] = 0;
disk_mem[17812] = 0;
disk_mem[17813] = 0;
disk_mem[17814] = 0;
disk_mem[17815] = 0;
disk_mem[17816] = 0;
disk_mem[17817] = 0;
disk_mem[17818] = 0;
disk_mem[17819] = 0;
disk_mem[17820] = 0;
disk_mem[17821] = 0;
disk_mem[17822] = 0;
disk_mem[17823] = 0;
disk_mem[17824] = 0;
disk_mem[17825] = 0;
disk_mem[17826] = 0;
disk_mem[17827] = 0;
disk_mem[17828] = 0;
disk_mem[17829] = 0;
disk_mem[17830] = 0;
disk_mem[17831] = 0;
disk_mem[17832] = 0;
disk_mem[17833] = 0;
disk_mem[17834] = 0;
disk_mem[17835] = 0;
disk_mem[17836] = 0;
disk_mem[17837] = 0;
disk_mem[17838] = 0;
disk_mem[17839] = 0;
disk_mem[17840] = 0;
disk_mem[17841] = 0;
disk_mem[17842] = 0;
disk_mem[17843] = 0;
disk_mem[17844] = 0;
disk_mem[17845] = 0;
disk_mem[17846] = 0;
disk_mem[17847] = 0;
disk_mem[17848] = 0;
disk_mem[17849] = 0;
disk_mem[17850] = 0;
disk_mem[17851] = 0;
disk_mem[17852] = 0;
disk_mem[17853] = 0;
disk_mem[17854] = 0;
disk_mem[17855] = 0;
disk_mem[17856] = 0;
disk_mem[17857] = 0;
disk_mem[17858] = 0;
disk_mem[17859] = 0;
disk_mem[17860] = 0;
disk_mem[17861] = 0;
disk_mem[17862] = 0;
disk_mem[17863] = 0;
disk_mem[17864] = 0;
disk_mem[17865] = 0;
disk_mem[17866] = 0;
disk_mem[17867] = 0;
disk_mem[17868] = 0;
disk_mem[17869] = 0;
disk_mem[17870] = 0;
disk_mem[17871] = 0;
disk_mem[17872] = 0;
disk_mem[17873] = 0;
disk_mem[17874] = 0;
disk_mem[17875] = 0;
disk_mem[17876] = 0;
disk_mem[17877] = 0;
disk_mem[17878] = 0;
disk_mem[17879] = 0;
disk_mem[17880] = 0;
disk_mem[17881] = 0;
disk_mem[17882] = 0;
disk_mem[17883] = 0;
disk_mem[17884] = 0;
disk_mem[17885] = 0;
disk_mem[17886] = 0;
disk_mem[17887] = 0;
disk_mem[17888] = 0;
disk_mem[17889] = 0;
disk_mem[17890] = 0;
disk_mem[17891] = 0;
disk_mem[17892] = 0;
disk_mem[17893] = 0;
disk_mem[17894] = 0;
disk_mem[17895] = 0;
disk_mem[17896] = 0;
disk_mem[17897] = 0;
disk_mem[17898] = 0;
disk_mem[17899] = 0;
disk_mem[17900] = 0;
disk_mem[17901] = 0;
disk_mem[17902] = 0;
disk_mem[17903] = 0;
disk_mem[17904] = 0;
disk_mem[17905] = 0;
disk_mem[17906] = 0;
disk_mem[17907] = 0;
disk_mem[17908] = 0;
disk_mem[17909] = 0;
disk_mem[17910] = 0;
disk_mem[17911] = 0;
disk_mem[17912] = 0;
disk_mem[17913] = 0;
disk_mem[17914] = 0;
disk_mem[17915] = 0;
disk_mem[17916] = 0;
disk_mem[17917] = 0;
disk_mem[17918] = 0;
disk_mem[17919] = 0;
disk_mem[17920] = 0;
disk_mem[17921] = 0;
disk_mem[17922] = 0;
disk_mem[17923] = 0;
disk_mem[17924] = 0;
disk_mem[17925] = 0;
disk_mem[17926] = 0;
disk_mem[17927] = 0;
disk_mem[17928] = 0;
disk_mem[17929] = 0;
disk_mem[17930] = 0;
disk_mem[17931] = 0;
disk_mem[17932] = 0;
disk_mem[17933] = 0;
disk_mem[17934] = 0;
disk_mem[17935] = 0;
disk_mem[17936] = 0;
disk_mem[17937] = 0;
disk_mem[17938] = 0;
disk_mem[17939] = 0;
disk_mem[17940] = 0;
disk_mem[17941] = 0;
disk_mem[17942] = 0;
disk_mem[17943] = 0;
disk_mem[17944] = 0;
disk_mem[17945] = 0;
disk_mem[17946] = 0;
disk_mem[17947] = 0;
disk_mem[17948] = 0;
disk_mem[17949] = 0;
disk_mem[17950] = 0;
disk_mem[17951] = 0;
disk_mem[17952] = 0;
disk_mem[17953] = 0;
disk_mem[17954] = 0;
disk_mem[17955] = 0;
disk_mem[17956] = 0;
disk_mem[17957] = 0;
disk_mem[17958] = 0;
disk_mem[17959] = 0;
disk_mem[17960] = 0;
disk_mem[17961] = 0;
disk_mem[17962] = 0;
disk_mem[17963] = 0;
disk_mem[17964] = 0;
disk_mem[17965] = 0;
disk_mem[17966] = 0;
disk_mem[17967] = 0;
disk_mem[17968] = 0;
disk_mem[17969] = 0;
disk_mem[17970] = 0;
disk_mem[17971] = 0;
disk_mem[17972] = 0;
disk_mem[17973] = 0;
disk_mem[17974] = 0;
disk_mem[17975] = 0;
disk_mem[17976] = 0;
disk_mem[17977] = 0;
disk_mem[17978] = 0;
disk_mem[17979] = 0;
disk_mem[17980] = 0;
disk_mem[17981] = 0;
disk_mem[17982] = 0;
disk_mem[17983] = 0;
disk_mem[17984] = 0;
disk_mem[17985] = 0;
disk_mem[17986] = 0;
disk_mem[17987] = 0;
disk_mem[17988] = 0;
disk_mem[17989] = 0;
disk_mem[17990] = 0;
disk_mem[17991] = 0;
disk_mem[17992] = 0;
disk_mem[17993] = 0;
disk_mem[17994] = 0;
disk_mem[17995] = 0;
disk_mem[17996] = 0;
disk_mem[17997] = 0;
disk_mem[17998] = 0;
disk_mem[17999] = 0;
disk_mem[18000] = 0;
disk_mem[18001] = 0;
disk_mem[18002] = 0;
disk_mem[18003] = 0;
disk_mem[18004] = 0;
disk_mem[18005] = 0;
disk_mem[18006] = 0;
disk_mem[18007] = 0;
disk_mem[18008] = 0;
disk_mem[18009] = 0;
disk_mem[18010] = 0;
disk_mem[18011] = 0;
disk_mem[18012] = 0;
disk_mem[18013] = 0;
disk_mem[18014] = 0;
disk_mem[18015] = 0;
disk_mem[18016] = 0;
disk_mem[18017] = 0;
disk_mem[18018] = 0;
disk_mem[18019] = 0;
disk_mem[18020] = 0;
disk_mem[18021] = 0;
disk_mem[18022] = 0;
disk_mem[18023] = 0;
disk_mem[18024] = 0;
disk_mem[18025] = 0;
disk_mem[18026] = 0;
disk_mem[18027] = 0;
disk_mem[18028] = 0;
disk_mem[18029] = 0;
disk_mem[18030] = 0;
disk_mem[18031] = 0;
disk_mem[18032] = 0;
disk_mem[18033] = 0;
disk_mem[18034] = 0;
disk_mem[18035] = 0;
disk_mem[18036] = 0;
disk_mem[18037] = 0;
disk_mem[18038] = 0;
disk_mem[18039] = 0;
disk_mem[18040] = 0;
disk_mem[18041] = 0;
disk_mem[18042] = 0;
disk_mem[18043] = 0;
disk_mem[18044] = 0;
disk_mem[18045] = 0;
disk_mem[18046] = 0;
disk_mem[18047] = 0;
disk_mem[18048] = 0;
disk_mem[18049] = 0;
disk_mem[18050] = 0;
disk_mem[18051] = 0;
disk_mem[18052] = 0;
disk_mem[18053] = 0;
disk_mem[18054] = 0;
disk_mem[18055] = 0;
disk_mem[18056] = 0;
disk_mem[18057] = 0;
disk_mem[18058] = 0;
disk_mem[18059] = 0;
disk_mem[18060] = 0;
disk_mem[18061] = 0;
disk_mem[18062] = 0;
disk_mem[18063] = 0;
disk_mem[18064] = 0;
disk_mem[18065] = 0;
disk_mem[18066] = 0;
disk_mem[18067] = 0;
disk_mem[18068] = 0;
disk_mem[18069] = 0;
disk_mem[18070] = 0;
disk_mem[18071] = 0;
disk_mem[18072] = 0;
disk_mem[18073] = 0;
disk_mem[18074] = 0;
disk_mem[18075] = 0;
disk_mem[18076] = 0;
disk_mem[18077] = 0;
disk_mem[18078] = 0;
disk_mem[18079] = 0;
disk_mem[18080] = 0;
disk_mem[18081] = 0;
disk_mem[18082] = 0;
disk_mem[18083] = 0;
disk_mem[18084] = 0;
disk_mem[18085] = 0;
disk_mem[18086] = 0;
disk_mem[18087] = 0;
disk_mem[18088] = 0;
disk_mem[18089] = 0;
disk_mem[18090] = 0;
disk_mem[18091] = 0;
disk_mem[18092] = 0;
disk_mem[18093] = 0;
disk_mem[18094] = 0;
disk_mem[18095] = 0;
disk_mem[18096] = 0;
disk_mem[18097] = 0;
disk_mem[18098] = 0;
disk_mem[18099] = 0;
disk_mem[18100] = 0;
disk_mem[18101] = 0;
disk_mem[18102] = 0;
disk_mem[18103] = 0;
disk_mem[18104] = 0;
disk_mem[18105] = 0;
disk_mem[18106] = 0;
disk_mem[18107] = 0;
disk_mem[18108] = 0;
disk_mem[18109] = 0;
disk_mem[18110] = 0;
disk_mem[18111] = 0;
disk_mem[18112] = 0;
disk_mem[18113] = 0;
disk_mem[18114] = 0;
disk_mem[18115] = 0;
disk_mem[18116] = 0;
disk_mem[18117] = 0;
disk_mem[18118] = 0;
disk_mem[18119] = 0;
disk_mem[18120] = 0;
disk_mem[18121] = 0;
disk_mem[18122] = 0;
disk_mem[18123] = 0;
disk_mem[18124] = 0;
disk_mem[18125] = 0;
disk_mem[18126] = 0;
disk_mem[18127] = 0;
disk_mem[18128] = 0;
disk_mem[18129] = 0;
disk_mem[18130] = 0;
disk_mem[18131] = 0;
disk_mem[18132] = 0;
disk_mem[18133] = 0;
disk_mem[18134] = 0;
disk_mem[18135] = 0;
disk_mem[18136] = 0;
disk_mem[18137] = 0;
disk_mem[18138] = 0;
disk_mem[18139] = 0;
disk_mem[18140] = 0;
disk_mem[18141] = 0;
disk_mem[18142] = 0;
disk_mem[18143] = 0;
disk_mem[18144] = 0;
disk_mem[18145] = 0;
disk_mem[18146] = 0;
disk_mem[18147] = 0;
disk_mem[18148] = 0;
disk_mem[18149] = 0;
disk_mem[18150] = 0;
disk_mem[18151] = 0;
disk_mem[18152] = 0;
disk_mem[18153] = 0;
disk_mem[18154] = 0;
disk_mem[18155] = 0;
disk_mem[18156] = 0;
disk_mem[18157] = 0;
disk_mem[18158] = 0;
disk_mem[18159] = 0;
disk_mem[18160] = 0;
disk_mem[18161] = 0;
disk_mem[18162] = 0;
disk_mem[18163] = 0;
disk_mem[18164] = 0;
disk_mem[18165] = 0;
disk_mem[18166] = 0;
disk_mem[18167] = 0;
disk_mem[18168] = 0;
disk_mem[18169] = 0;
disk_mem[18170] = 0;
disk_mem[18171] = 0;
disk_mem[18172] = 0;
disk_mem[18173] = 0;
disk_mem[18174] = 0;
disk_mem[18175] = 0;
disk_mem[18176] = 0;
disk_mem[18177] = 0;
disk_mem[18178] = 0;
disk_mem[18179] = 0;
disk_mem[18180] = 0;
disk_mem[18181] = 0;
disk_mem[18182] = 0;
disk_mem[18183] = 0;
disk_mem[18184] = 0;
disk_mem[18185] = 0;
disk_mem[18186] = 0;
disk_mem[18187] = 0;
disk_mem[18188] = 0;
disk_mem[18189] = 0;
disk_mem[18190] = 0;
disk_mem[18191] = 0;
disk_mem[18192] = 0;
disk_mem[18193] = 0;
disk_mem[18194] = 0;
disk_mem[18195] = 0;
disk_mem[18196] = 0;
disk_mem[18197] = 0;
disk_mem[18198] = 0;
disk_mem[18199] = 0;
disk_mem[18200] = 0;
disk_mem[18201] = 0;
disk_mem[18202] = 0;
disk_mem[18203] = 0;
disk_mem[18204] = 0;
disk_mem[18205] = 0;
disk_mem[18206] = 0;
disk_mem[18207] = 0;
disk_mem[18208] = 0;
disk_mem[18209] = 0;
disk_mem[18210] = 0;
disk_mem[18211] = 0;
disk_mem[18212] = 0;
disk_mem[18213] = 0;
disk_mem[18214] = 0;
disk_mem[18215] = 0;
disk_mem[18216] = 0;
disk_mem[18217] = 0;
disk_mem[18218] = 0;
disk_mem[18219] = 0;
disk_mem[18220] = 0;
disk_mem[18221] = 0;
disk_mem[18222] = 0;
disk_mem[18223] = 0;
disk_mem[18224] = 0;
disk_mem[18225] = 0;
disk_mem[18226] = 0;
disk_mem[18227] = 0;
disk_mem[18228] = 0;
disk_mem[18229] = 0;
disk_mem[18230] = 0;
disk_mem[18231] = 0;
disk_mem[18232] = 0;
disk_mem[18233] = 0;
disk_mem[18234] = 0;
disk_mem[18235] = 0;
disk_mem[18236] = 0;
disk_mem[18237] = 0;
disk_mem[18238] = 0;
disk_mem[18239] = 0;
disk_mem[18240] = 0;
disk_mem[18241] = 0;
disk_mem[18242] = 0;
disk_mem[18243] = 0;
disk_mem[18244] = 0;
disk_mem[18245] = 0;
disk_mem[18246] = 0;
disk_mem[18247] = 0;
disk_mem[18248] = 0;
disk_mem[18249] = 0;
disk_mem[18250] = 0;
disk_mem[18251] = 0;
disk_mem[18252] = 0;
disk_mem[18253] = 0;
disk_mem[18254] = 0;
disk_mem[18255] = 0;
disk_mem[18256] = 0;
disk_mem[18257] = 0;
disk_mem[18258] = 0;
disk_mem[18259] = 0;
disk_mem[18260] = 0;
disk_mem[18261] = 0;
disk_mem[18262] = 0;
disk_mem[18263] = 0;
disk_mem[18264] = 0;
disk_mem[18265] = 0;
disk_mem[18266] = 0;
disk_mem[18267] = 0;
disk_mem[18268] = 0;
disk_mem[18269] = 0;
disk_mem[18270] = 0;
disk_mem[18271] = 0;
disk_mem[18272] = 0;
disk_mem[18273] = 0;
disk_mem[18274] = 0;
disk_mem[18275] = 0;
disk_mem[18276] = 0;
disk_mem[18277] = 0;
disk_mem[18278] = 0;
disk_mem[18279] = 0;
disk_mem[18280] = 0;
disk_mem[18281] = 0;
disk_mem[18282] = 0;
disk_mem[18283] = 0;
disk_mem[18284] = 0;
disk_mem[18285] = 0;
disk_mem[18286] = 0;
disk_mem[18287] = 0;
disk_mem[18288] = 0;
disk_mem[18289] = 0;
disk_mem[18290] = 0;
disk_mem[18291] = 0;
disk_mem[18292] = 0;
disk_mem[18293] = 0;
disk_mem[18294] = 0;
disk_mem[18295] = 0;
disk_mem[18296] = 0;
disk_mem[18297] = 0;
disk_mem[18298] = 0;
disk_mem[18299] = 0;
disk_mem[18300] = 0;
disk_mem[18301] = 0;
disk_mem[18302] = 0;
disk_mem[18303] = 0;
disk_mem[18304] = 0;
disk_mem[18305] = 0;
disk_mem[18306] = 0;
disk_mem[18307] = 0;
disk_mem[18308] = 0;
disk_mem[18309] = 0;
disk_mem[18310] = 0;
disk_mem[18311] = 0;
disk_mem[18312] = 0;
disk_mem[18313] = 0;
disk_mem[18314] = 0;
disk_mem[18315] = 0;
disk_mem[18316] = 0;
disk_mem[18317] = 0;
disk_mem[18318] = 0;
disk_mem[18319] = 0;
disk_mem[18320] = 0;
disk_mem[18321] = 0;
disk_mem[18322] = 0;
disk_mem[18323] = 0;
disk_mem[18324] = 0;
disk_mem[18325] = 0;
disk_mem[18326] = 0;
disk_mem[18327] = 0;
disk_mem[18328] = 0;
disk_mem[18329] = 0;
disk_mem[18330] = 0;
disk_mem[18331] = 0;
disk_mem[18332] = 0;
disk_mem[18333] = 0;
disk_mem[18334] = 0;
disk_mem[18335] = 0;
disk_mem[18336] = 0;
disk_mem[18337] = 0;
disk_mem[18338] = 0;
disk_mem[18339] = 0;
disk_mem[18340] = 0;
disk_mem[18341] = 0;
disk_mem[18342] = 0;
disk_mem[18343] = 0;
disk_mem[18344] = 0;
disk_mem[18345] = 0;
disk_mem[18346] = 0;
disk_mem[18347] = 0;
disk_mem[18348] = 0;
disk_mem[18349] = 0;
disk_mem[18350] = 0;
disk_mem[18351] = 0;
disk_mem[18352] = 0;
disk_mem[18353] = 0;
disk_mem[18354] = 0;
disk_mem[18355] = 0;
disk_mem[18356] = 0;
disk_mem[18357] = 0;
disk_mem[18358] = 0;
disk_mem[18359] = 0;
disk_mem[18360] = 0;
disk_mem[18361] = 0;
disk_mem[18362] = 0;
disk_mem[18363] = 0;
disk_mem[18364] = 0;
disk_mem[18365] = 0;
disk_mem[18366] = 0;
disk_mem[18367] = 0;
disk_mem[18368] = 0;
disk_mem[18369] = 0;
disk_mem[18370] = 0;
disk_mem[18371] = 0;
disk_mem[18372] = 0;
disk_mem[18373] = 0;
disk_mem[18374] = 0;
disk_mem[18375] = 0;
disk_mem[18376] = 0;
disk_mem[18377] = 0;
disk_mem[18378] = 0;
disk_mem[18379] = 0;
disk_mem[18380] = 0;
disk_mem[18381] = 0;
disk_mem[18382] = 0;
disk_mem[18383] = 0;
disk_mem[18384] = 0;
disk_mem[18385] = 0;
disk_mem[18386] = 0;
disk_mem[18387] = 0;
disk_mem[18388] = 0;
disk_mem[18389] = 0;
disk_mem[18390] = 0;
disk_mem[18391] = 0;
disk_mem[18392] = 0;
disk_mem[18393] = 0;
disk_mem[18394] = 0;
disk_mem[18395] = 0;
disk_mem[18396] = 0;
disk_mem[18397] = 0;
disk_mem[18398] = 0;
disk_mem[18399] = 0;
disk_mem[18400] = 0;
disk_mem[18401] = 0;
disk_mem[18402] = 0;
disk_mem[18403] = 0;
disk_mem[18404] = 0;
disk_mem[18405] = 0;
disk_mem[18406] = 0;
disk_mem[18407] = 0;
disk_mem[18408] = 0;
disk_mem[18409] = 0;
disk_mem[18410] = 0;
disk_mem[18411] = 0;
disk_mem[18412] = 0;
disk_mem[18413] = 0;
disk_mem[18414] = 0;
disk_mem[18415] = 0;
disk_mem[18416] = 0;
disk_mem[18417] = 0;
disk_mem[18418] = 0;
disk_mem[18419] = 0;
disk_mem[18420] = 0;
disk_mem[18421] = 0;
disk_mem[18422] = 0;
disk_mem[18423] = 0;
disk_mem[18424] = 0;
disk_mem[18425] = 0;
disk_mem[18426] = 0;
disk_mem[18427] = 0;
disk_mem[18428] = 0;
disk_mem[18429] = 0;
disk_mem[18430] = 0;
disk_mem[18431] = 0;
disk_mem[18432] = 0;
disk_mem[18433] = 0;
disk_mem[18434] = 0;
disk_mem[18435] = 0;
disk_mem[18436] = 0;
disk_mem[18437] = 0;
disk_mem[18438] = 0;
disk_mem[18439] = 0;
disk_mem[18440] = 0;
disk_mem[18441] = 0;
disk_mem[18442] = 0;
disk_mem[18443] = 0;
disk_mem[18444] = 0;
disk_mem[18445] = 0;
disk_mem[18446] = 0;
disk_mem[18447] = 0;
disk_mem[18448] = 0;
disk_mem[18449] = 0;
disk_mem[18450] = 0;
disk_mem[18451] = 0;
disk_mem[18452] = 0;
disk_mem[18453] = 0;
disk_mem[18454] = 0;
disk_mem[18455] = 0;
disk_mem[18456] = 0;
disk_mem[18457] = 0;
disk_mem[18458] = 0;
disk_mem[18459] = 0;
disk_mem[18460] = 0;
disk_mem[18461] = 0;
disk_mem[18462] = 0;
disk_mem[18463] = 0;
disk_mem[18464] = 0;
disk_mem[18465] = 0;
disk_mem[18466] = 0;
disk_mem[18467] = 0;
disk_mem[18468] = 0;
disk_mem[18469] = 0;
disk_mem[18470] = 0;
disk_mem[18471] = 0;
disk_mem[18472] = 0;
disk_mem[18473] = 0;
disk_mem[18474] = 0;
disk_mem[18475] = 0;
disk_mem[18476] = 0;
disk_mem[18477] = 0;
disk_mem[18478] = 0;
disk_mem[18479] = 0;
disk_mem[18480] = 0;
disk_mem[18481] = 0;
disk_mem[18482] = 0;
disk_mem[18483] = 0;
disk_mem[18484] = 0;
disk_mem[18485] = 0;
disk_mem[18486] = 0;
disk_mem[18487] = 0;
disk_mem[18488] = 0;
disk_mem[18489] = 0;
disk_mem[18490] = 0;
disk_mem[18491] = 0;
disk_mem[18492] = 0;
disk_mem[18493] = 0;
disk_mem[18494] = 0;
disk_mem[18495] = 0;
disk_mem[18496] = 0;
disk_mem[18497] = 0;
disk_mem[18498] = 0;
disk_mem[18499] = 0;
disk_mem[18500] = 0;
disk_mem[18501] = 0;
disk_mem[18502] = 0;
disk_mem[18503] = 0;
disk_mem[18504] = 0;
disk_mem[18505] = 0;
disk_mem[18506] = 0;
disk_mem[18507] = 0;
disk_mem[18508] = 0;
disk_mem[18509] = 0;
disk_mem[18510] = 0;
disk_mem[18511] = 0;
disk_mem[18512] = 0;
disk_mem[18513] = 0;
disk_mem[18514] = 0;
disk_mem[18515] = 0;
disk_mem[18516] = 0;
disk_mem[18517] = 0;
disk_mem[18518] = 0;
disk_mem[18519] = 0;
disk_mem[18520] = 0;
disk_mem[18521] = 0;
disk_mem[18522] = 0;
disk_mem[18523] = 0;
disk_mem[18524] = 0;
disk_mem[18525] = 0;
disk_mem[18526] = 0;
disk_mem[18527] = 0;
disk_mem[18528] = 0;
disk_mem[18529] = 0;
disk_mem[18530] = 0;
disk_mem[18531] = 0;
disk_mem[18532] = 0;
disk_mem[18533] = 0;
disk_mem[18534] = 0;
disk_mem[18535] = 0;
disk_mem[18536] = 0;
disk_mem[18537] = 0;
disk_mem[18538] = 0;
disk_mem[18539] = 0;
disk_mem[18540] = 0;
disk_mem[18541] = 0;
disk_mem[18542] = 0;
disk_mem[18543] = 0;
disk_mem[18544] = 0;
disk_mem[18545] = 0;
disk_mem[18546] = 0;
disk_mem[18547] = 0;
disk_mem[18548] = 0;
disk_mem[18549] = 0;
disk_mem[18550] = 0;
disk_mem[18551] = 0;
disk_mem[18552] = 0;
disk_mem[18553] = 0;
disk_mem[18554] = 0;
disk_mem[18555] = 0;
disk_mem[18556] = 0;
disk_mem[18557] = 0;
disk_mem[18558] = 0;
disk_mem[18559] = 0;
disk_mem[18560] = 0;
disk_mem[18561] = 0;
disk_mem[18562] = 0;
disk_mem[18563] = 0;
disk_mem[18564] = 0;
disk_mem[18565] = 0;
disk_mem[18566] = 0;
disk_mem[18567] = 0;
disk_mem[18568] = 0;
disk_mem[18569] = 0;
disk_mem[18570] = 0;
disk_mem[18571] = 0;
disk_mem[18572] = 0;
disk_mem[18573] = 0;
disk_mem[18574] = 0;
disk_mem[18575] = 0;
disk_mem[18576] = 0;
disk_mem[18577] = 0;
disk_mem[18578] = 0;
disk_mem[18579] = 0;
disk_mem[18580] = 0;
disk_mem[18581] = 0;
disk_mem[18582] = 0;
disk_mem[18583] = 0;
disk_mem[18584] = 0;
disk_mem[18585] = 0;
disk_mem[18586] = 0;
disk_mem[18587] = 0;
disk_mem[18588] = 0;
disk_mem[18589] = 0;
disk_mem[18590] = 0;
disk_mem[18591] = 0;
disk_mem[18592] = 0;
disk_mem[18593] = 0;
disk_mem[18594] = 0;
disk_mem[18595] = 0;
disk_mem[18596] = 0;
disk_mem[18597] = 0;
disk_mem[18598] = 0;
disk_mem[18599] = 0;
disk_mem[18600] = 0;
disk_mem[18601] = 0;
disk_mem[18602] = 0;
disk_mem[18603] = 0;
disk_mem[18604] = 0;
disk_mem[18605] = 0;
disk_mem[18606] = 0;
disk_mem[18607] = 0;
disk_mem[18608] = 0;
disk_mem[18609] = 0;
disk_mem[18610] = 0;
disk_mem[18611] = 0;
disk_mem[18612] = 0;
disk_mem[18613] = 0;
disk_mem[18614] = 0;
disk_mem[18615] = 0;
disk_mem[18616] = 0;
disk_mem[18617] = 0;
disk_mem[18618] = 0;
disk_mem[18619] = 0;
disk_mem[18620] = 0;
disk_mem[18621] = 0;
disk_mem[18622] = 0;
disk_mem[18623] = 0;
disk_mem[18624] = 0;
disk_mem[18625] = 0;
disk_mem[18626] = 0;
disk_mem[18627] = 0;
disk_mem[18628] = 0;
disk_mem[18629] = 0;
disk_mem[18630] = 0;
disk_mem[18631] = 0;
disk_mem[18632] = 0;
disk_mem[18633] = 0;
disk_mem[18634] = 0;
disk_mem[18635] = 0;
disk_mem[18636] = 0;
disk_mem[18637] = 0;
disk_mem[18638] = 0;
disk_mem[18639] = 0;
disk_mem[18640] = 0;
disk_mem[18641] = 0;
disk_mem[18642] = 0;
disk_mem[18643] = 0;
disk_mem[18644] = 0;
disk_mem[18645] = 0;
disk_mem[18646] = 0;
disk_mem[18647] = 0;
disk_mem[18648] = 0;
disk_mem[18649] = 0;
disk_mem[18650] = 0;
disk_mem[18651] = 0;
disk_mem[18652] = 0;
disk_mem[18653] = 0;
disk_mem[18654] = 0;
disk_mem[18655] = 0;
disk_mem[18656] = 0;
disk_mem[18657] = 0;
disk_mem[18658] = 0;
disk_mem[18659] = 0;
disk_mem[18660] = 0;
disk_mem[18661] = 0;
disk_mem[18662] = 0;
disk_mem[18663] = 0;
disk_mem[18664] = 0;
disk_mem[18665] = 0;
disk_mem[18666] = 0;
disk_mem[18667] = 0;
disk_mem[18668] = 0;
disk_mem[18669] = 0;
disk_mem[18670] = 0;
disk_mem[18671] = 0;
disk_mem[18672] = 0;
disk_mem[18673] = 0;
disk_mem[18674] = 0;
disk_mem[18675] = 0;
disk_mem[18676] = 0;
disk_mem[18677] = 0;
disk_mem[18678] = 0;
disk_mem[18679] = 0;
disk_mem[18680] = 0;
disk_mem[18681] = 0;
disk_mem[18682] = 0;
disk_mem[18683] = 0;
disk_mem[18684] = 0;
disk_mem[18685] = 0;
disk_mem[18686] = 0;
disk_mem[18687] = 0;
disk_mem[18688] = 0;
disk_mem[18689] = 0;
disk_mem[18690] = 0;
disk_mem[18691] = 0;
disk_mem[18692] = 0;
disk_mem[18693] = 0;
disk_mem[18694] = 0;
disk_mem[18695] = 0;
disk_mem[18696] = 0;
disk_mem[18697] = 0;
disk_mem[18698] = 0;
disk_mem[18699] = 0;
disk_mem[18700] = 0;
disk_mem[18701] = 0;
disk_mem[18702] = 0;
disk_mem[18703] = 0;
disk_mem[18704] = 0;
disk_mem[18705] = 0;
disk_mem[18706] = 0;
disk_mem[18707] = 0;
disk_mem[18708] = 0;
disk_mem[18709] = 0;
disk_mem[18710] = 0;
disk_mem[18711] = 0;
disk_mem[18712] = 0;
disk_mem[18713] = 0;
disk_mem[18714] = 0;
disk_mem[18715] = 0;
disk_mem[18716] = 0;
disk_mem[18717] = 0;
disk_mem[18718] = 0;
disk_mem[18719] = 0;
disk_mem[18720] = 0;
disk_mem[18721] = 0;
disk_mem[18722] = 0;
disk_mem[18723] = 0;
disk_mem[18724] = 0;
disk_mem[18725] = 0;
disk_mem[18726] = 0;
disk_mem[18727] = 0;
disk_mem[18728] = 0;
disk_mem[18729] = 0;
disk_mem[18730] = 0;
disk_mem[18731] = 0;
disk_mem[18732] = 0;
disk_mem[18733] = 0;
disk_mem[18734] = 0;
disk_mem[18735] = 0;
disk_mem[18736] = 0;
disk_mem[18737] = 0;
disk_mem[18738] = 0;
disk_mem[18739] = 0;
disk_mem[18740] = 0;
disk_mem[18741] = 0;
disk_mem[18742] = 0;
disk_mem[18743] = 0;
disk_mem[18744] = 0;
disk_mem[18745] = 0;
disk_mem[18746] = 0;
disk_mem[18747] = 0;
disk_mem[18748] = 0;
disk_mem[18749] = 0;
disk_mem[18750] = 0;
disk_mem[18751] = 0;
disk_mem[18752] = 0;
disk_mem[18753] = 0;
disk_mem[18754] = 0;
disk_mem[18755] = 0;
disk_mem[18756] = 0;
disk_mem[18757] = 0;
disk_mem[18758] = 0;
disk_mem[18759] = 0;
disk_mem[18760] = 0;
disk_mem[18761] = 0;
disk_mem[18762] = 0;
disk_mem[18763] = 0;
disk_mem[18764] = 0;
disk_mem[18765] = 0;
disk_mem[18766] = 0;
disk_mem[18767] = 0;
disk_mem[18768] = 0;
disk_mem[18769] = 0;
disk_mem[18770] = 0;
disk_mem[18771] = 0;
disk_mem[18772] = 0;
disk_mem[18773] = 0;
disk_mem[18774] = 0;
disk_mem[18775] = 0;
disk_mem[18776] = 0;
disk_mem[18777] = 0;
disk_mem[18778] = 0;
disk_mem[18779] = 0;
disk_mem[18780] = 0;
disk_mem[18781] = 0;
disk_mem[18782] = 0;
disk_mem[18783] = 0;
disk_mem[18784] = 0;
disk_mem[18785] = 0;
disk_mem[18786] = 0;
disk_mem[18787] = 0;
disk_mem[18788] = 0;
disk_mem[18789] = 0;
disk_mem[18790] = 0;
disk_mem[18791] = 0;
disk_mem[18792] = 0;
disk_mem[18793] = 0;
disk_mem[18794] = 0;
disk_mem[18795] = 0;
disk_mem[18796] = 0;
disk_mem[18797] = 0;
disk_mem[18798] = 0;
disk_mem[18799] = 0;
disk_mem[18800] = 0;
disk_mem[18801] = 0;
disk_mem[18802] = 0;
disk_mem[18803] = 0;
disk_mem[18804] = 0;
disk_mem[18805] = 0;
disk_mem[18806] = 0;
disk_mem[18807] = 0;
disk_mem[18808] = 0;
disk_mem[18809] = 0;
disk_mem[18810] = 0;
disk_mem[18811] = 0;
disk_mem[18812] = 0;
disk_mem[18813] = 0;
disk_mem[18814] = 0;
disk_mem[18815] = 0;
disk_mem[18816] = 0;
disk_mem[18817] = 0;
disk_mem[18818] = 0;
disk_mem[18819] = 0;
disk_mem[18820] = 0;
disk_mem[18821] = 0;
disk_mem[18822] = 0;
disk_mem[18823] = 0;
disk_mem[18824] = 0;
disk_mem[18825] = 0;
disk_mem[18826] = 0;
disk_mem[18827] = 0;
disk_mem[18828] = 0;
disk_mem[18829] = 0;
disk_mem[18830] = 0;
disk_mem[18831] = 0;
disk_mem[18832] = 0;
disk_mem[18833] = 0;
disk_mem[18834] = 0;
disk_mem[18835] = 0;
disk_mem[18836] = 0;
disk_mem[18837] = 0;
disk_mem[18838] = 0;
disk_mem[18839] = 0;
disk_mem[18840] = 0;
disk_mem[18841] = 0;
disk_mem[18842] = 0;
disk_mem[18843] = 0;
disk_mem[18844] = 0;
disk_mem[18845] = 0;
disk_mem[18846] = 0;
disk_mem[18847] = 0;
disk_mem[18848] = 0;
disk_mem[18849] = 0;
disk_mem[18850] = 0;
disk_mem[18851] = 0;
disk_mem[18852] = 0;
disk_mem[18853] = 0;
disk_mem[18854] = 0;
disk_mem[18855] = 0;
disk_mem[18856] = 0;
disk_mem[18857] = 0;
disk_mem[18858] = 0;
disk_mem[18859] = 0;
disk_mem[18860] = 0;
disk_mem[18861] = 0;
disk_mem[18862] = 0;
disk_mem[18863] = 0;
disk_mem[18864] = 0;
disk_mem[18865] = 0;
disk_mem[18866] = 0;
disk_mem[18867] = 0;
disk_mem[18868] = 0;
disk_mem[18869] = 0;
disk_mem[18870] = 0;
disk_mem[18871] = 0;
disk_mem[18872] = 0;
disk_mem[18873] = 0;
disk_mem[18874] = 0;
disk_mem[18875] = 0;
disk_mem[18876] = 0;
disk_mem[18877] = 0;
disk_mem[18878] = 0;
disk_mem[18879] = 0;
disk_mem[18880] = 0;
disk_mem[18881] = 0;
disk_mem[18882] = 0;
disk_mem[18883] = 0;
disk_mem[18884] = 0;
disk_mem[18885] = 0;
disk_mem[18886] = 0;
disk_mem[18887] = 0;
disk_mem[18888] = 0;
disk_mem[18889] = 0;
disk_mem[18890] = 0;
disk_mem[18891] = 0;
disk_mem[18892] = 0;
disk_mem[18893] = 0;
disk_mem[18894] = 0;
disk_mem[18895] = 0;
disk_mem[18896] = 0;
disk_mem[18897] = 0;
disk_mem[18898] = 0;
disk_mem[18899] = 0;
disk_mem[18900] = 0;
disk_mem[18901] = 0;
disk_mem[18902] = 0;
disk_mem[18903] = 0;
disk_mem[18904] = 0;
disk_mem[18905] = 0;
disk_mem[18906] = 0;
disk_mem[18907] = 0;
disk_mem[18908] = 0;
disk_mem[18909] = 0;
disk_mem[18910] = 0;
disk_mem[18911] = 0;
disk_mem[18912] = 0;
disk_mem[18913] = 0;
disk_mem[18914] = 0;
disk_mem[18915] = 0;
disk_mem[18916] = 0;
disk_mem[18917] = 0;
disk_mem[18918] = 0;
disk_mem[18919] = 0;
disk_mem[18920] = 0;
disk_mem[18921] = 0;
disk_mem[18922] = 0;
disk_mem[18923] = 0;
disk_mem[18924] = 0;
disk_mem[18925] = 0;
disk_mem[18926] = 0;
disk_mem[18927] = 0;
disk_mem[18928] = 0;
disk_mem[18929] = 0;
disk_mem[18930] = 0;
disk_mem[18931] = 0;
disk_mem[18932] = 0;
disk_mem[18933] = 0;
disk_mem[18934] = 0;
disk_mem[18935] = 0;
disk_mem[18936] = 0;
disk_mem[18937] = 0;
disk_mem[18938] = 0;
disk_mem[18939] = 0;
disk_mem[18940] = 0;
disk_mem[18941] = 0;
disk_mem[18942] = 0;
disk_mem[18943] = 0;
disk_mem[18944] = 0;
disk_mem[18945] = 0;
disk_mem[18946] = 0;
disk_mem[18947] = 0;
disk_mem[18948] = 0;
disk_mem[18949] = 0;
disk_mem[18950] = 0;
disk_mem[18951] = 0;
disk_mem[18952] = 0;
disk_mem[18953] = 0;
disk_mem[18954] = 0;
disk_mem[18955] = 0;
disk_mem[18956] = 0;
disk_mem[18957] = 0;
disk_mem[18958] = 0;
disk_mem[18959] = 0;
disk_mem[18960] = 0;
disk_mem[18961] = 0;
disk_mem[18962] = 0;
disk_mem[18963] = 0;
disk_mem[18964] = 0;
disk_mem[18965] = 0;
disk_mem[18966] = 0;
disk_mem[18967] = 0;
disk_mem[18968] = 0;
disk_mem[18969] = 0;
disk_mem[18970] = 0;
disk_mem[18971] = 0;
disk_mem[18972] = 0;
disk_mem[18973] = 0;
disk_mem[18974] = 0;
disk_mem[18975] = 0;
disk_mem[18976] = 0;
disk_mem[18977] = 0;
disk_mem[18978] = 0;
disk_mem[18979] = 0;
disk_mem[18980] = 0;
disk_mem[18981] = 0;
disk_mem[18982] = 0;
disk_mem[18983] = 0;
disk_mem[18984] = 0;
disk_mem[18985] = 0;
disk_mem[18986] = 0;
disk_mem[18987] = 0;
disk_mem[18988] = 0;
disk_mem[18989] = 0;
disk_mem[18990] = 0;
disk_mem[18991] = 0;
disk_mem[18992] = 0;
disk_mem[18993] = 0;
disk_mem[18994] = 0;
disk_mem[18995] = 0;
disk_mem[18996] = 0;
disk_mem[18997] = 0;
disk_mem[18998] = 0;
disk_mem[18999] = 0;
disk_mem[19000] = 0;
disk_mem[19001] = 0;
disk_mem[19002] = 0;
disk_mem[19003] = 0;
disk_mem[19004] = 0;
disk_mem[19005] = 0;
disk_mem[19006] = 0;
disk_mem[19007] = 0;
disk_mem[19008] = 0;
disk_mem[19009] = 0;
disk_mem[19010] = 0;
disk_mem[19011] = 0;
disk_mem[19012] = 0;
disk_mem[19013] = 0;
disk_mem[19014] = 0;
disk_mem[19015] = 0;
disk_mem[19016] = 0;
disk_mem[19017] = 0;
disk_mem[19018] = 0;
disk_mem[19019] = 0;
disk_mem[19020] = 0;
disk_mem[19021] = 0;
disk_mem[19022] = 0;
disk_mem[19023] = 0;
disk_mem[19024] = 0;
disk_mem[19025] = 0;
disk_mem[19026] = 0;
disk_mem[19027] = 0;
disk_mem[19028] = 0;
disk_mem[19029] = 0;
disk_mem[19030] = 0;
disk_mem[19031] = 0;
disk_mem[19032] = 0;
disk_mem[19033] = 0;
disk_mem[19034] = 0;
disk_mem[19035] = 0;
disk_mem[19036] = 0;
disk_mem[19037] = 0;
disk_mem[19038] = 0;
disk_mem[19039] = 0;
disk_mem[19040] = 0;
disk_mem[19041] = 0;
disk_mem[19042] = 0;
disk_mem[19043] = 0;
disk_mem[19044] = 0;
disk_mem[19045] = 0;
disk_mem[19046] = 0;
disk_mem[19047] = 0;
disk_mem[19048] = 0;
disk_mem[19049] = 0;
disk_mem[19050] = 0;
disk_mem[19051] = 0;
disk_mem[19052] = 0;
disk_mem[19053] = 0;
disk_mem[19054] = 0;
disk_mem[19055] = 0;
disk_mem[19056] = 0;
disk_mem[19057] = 0;
disk_mem[19058] = 0;
disk_mem[19059] = 0;
disk_mem[19060] = 0;
disk_mem[19061] = 0;
disk_mem[19062] = 0;
disk_mem[19063] = 0;
disk_mem[19064] = 0;
disk_mem[19065] = 0;
disk_mem[19066] = 0;
disk_mem[19067] = 0;
disk_mem[19068] = 0;
disk_mem[19069] = 0;
disk_mem[19070] = 0;
disk_mem[19071] = 0;
disk_mem[19072] = 0;
disk_mem[19073] = 0;
disk_mem[19074] = 0;
disk_mem[19075] = 0;
disk_mem[19076] = 0;
disk_mem[19077] = 0;
disk_mem[19078] = 0;
disk_mem[19079] = 0;
disk_mem[19080] = 0;
disk_mem[19081] = 0;
disk_mem[19082] = 0;
disk_mem[19083] = 0;
disk_mem[19084] = 0;
disk_mem[19085] = 0;
disk_mem[19086] = 0;
disk_mem[19087] = 0;
disk_mem[19088] = 0;
disk_mem[19089] = 0;
disk_mem[19090] = 0;
disk_mem[19091] = 0;
disk_mem[19092] = 0;
disk_mem[19093] = 0;
disk_mem[19094] = 0;
disk_mem[19095] = 0;
disk_mem[19096] = 0;
disk_mem[19097] = 0;
disk_mem[19098] = 0;
disk_mem[19099] = 0;
disk_mem[19100] = 0;
disk_mem[19101] = 0;
disk_mem[19102] = 0;
disk_mem[19103] = 0;
disk_mem[19104] = 0;
disk_mem[19105] = 0;
disk_mem[19106] = 0;
disk_mem[19107] = 0;
disk_mem[19108] = 0;
disk_mem[19109] = 0;
disk_mem[19110] = 0;
disk_mem[19111] = 0;
disk_mem[19112] = 0;
disk_mem[19113] = 0;
disk_mem[19114] = 0;
disk_mem[19115] = 0;
disk_mem[19116] = 0;
disk_mem[19117] = 0;
disk_mem[19118] = 0;
disk_mem[19119] = 0;
disk_mem[19120] = 0;
disk_mem[19121] = 0;
disk_mem[19122] = 0;
disk_mem[19123] = 0;
disk_mem[19124] = 0;
disk_mem[19125] = 0;
disk_mem[19126] = 0;
disk_mem[19127] = 0;
disk_mem[19128] = 0;
disk_mem[19129] = 0;
disk_mem[19130] = 0;
disk_mem[19131] = 0;
disk_mem[19132] = 0;
disk_mem[19133] = 0;
disk_mem[19134] = 0;
disk_mem[19135] = 0;
disk_mem[19136] = 0;
disk_mem[19137] = 0;
disk_mem[19138] = 0;
disk_mem[19139] = 0;
disk_mem[19140] = 0;
disk_mem[19141] = 0;
disk_mem[19142] = 0;
disk_mem[19143] = 0;
disk_mem[19144] = 0;
disk_mem[19145] = 0;
disk_mem[19146] = 0;
disk_mem[19147] = 0;
disk_mem[19148] = 0;
disk_mem[19149] = 0;
disk_mem[19150] = 0;
disk_mem[19151] = 0;
disk_mem[19152] = 0;
disk_mem[19153] = 0;
disk_mem[19154] = 0;
disk_mem[19155] = 0;
disk_mem[19156] = 0;
disk_mem[19157] = 0;
disk_mem[19158] = 0;
disk_mem[19159] = 0;
disk_mem[19160] = 0;
disk_mem[19161] = 0;
disk_mem[19162] = 0;
disk_mem[19163] = 0;
disk_mem[19164] = 0;
disk_mem[19165] = 0;
disk_mem[19166] = 0;
disk_mem[19167] = 0;
disk_mem[19168] = 0;
disk_mem[19169] = 0;
disk_mem[19170] = 0;
disk_mem[19171] = 0;
disk_mem[19172] = 0;
disk_mem[19173] = 0;
disk_mem[19174] = 0;
disk_mem[19175] = 0;
disk_mem[19176] = 0;
disk_mem[19177] = 0;
disk_mem[19178] = 0;
disk_mem[19179] = 0;
disk_mem[19180] = 0;
disk_mem[19181] = 0;
disk_mem[19182] = 0;
disk_mem[19183] = 0;
disk_mem[19184] = 0;
disk_mem[19185] = 0;
disk_mem[19186] = 0;
disk_mem[19187] = 0;
disk_mem[19188] = 0;
disk_mem[19189] = 0;
disk_mem[19190] = 0;
disk_mem[19191] = 0;
disk_mem[19192] = 0;
disk_mem[19193] = 0;
disk_mem[19194] = 0;
disk_mem[19195] = 0;
disk_mem[19196] = 0;
disk_mem[19197] = 0;
disk_mem[19198] = 0;
disk_mem[19199] = 0;
disk_mem[19200] = 0;
disk_mem[19201] = 0;
disk_mem[19202] = 0;
disk_mem[19203] = 0;
disk_mem[19204] = 0;
disk_mem[19205] = 0;
disk_mem[19206] = 0;
disk_mem[19207] = 0;
disk_mem[19208] = 0;
disk_mem[19209] = 0;
disk_mem[19210] = 0;
disk_mem[19211] = 0;
disk_mem[19212] = 0;
disk_mem[19213] = 0;
disk_mem[19214] = 0;
disk_mem[19215] = 0;
disk_mem[19216] = 0;
disk_mem[19217] = 0;
disk_mem[19218] = 0;
disk_mem[19219] = 0;
disk_mem[19220] = 0;
disk_mem[19221] = 0;
disk_mem[19222] = 0;
disk_mem[19223] = 0;
disk_mem[19224] = 0;
disk_mem[19225] = 0;
disk_mem[19226] = 0;
disk_mem[19227] = 0;
disk_mem[19228] = 0;
disk_mem[19229] = 0;
disk_mem[19230] = 0;
disk_mem[19231] = 0;
disk_mem[19232] = 0;
disk_mem[19233] = 0;
disk_mem[19234] = 0;
disk_mem[19235] = 0;
disk_mem[19236] = 0;
disk_mem[19237] = 0;
disk_mem[19238] = 0;
disk_mem[19239] = 0;
disk_mem[19240] = 0;
disk_mem[19241] = 0;
disk_mem[19242] = 0;
disk_mem[19243] = 0;
disk_mem[19244] = 0;
disk_mem[19245] = 0;
disk_mem[19246] = 0;
disk_mem[19247] = 0;
disk_mem[19248] = 0;
disk_mem[19249] = 0;
disk_mem[19250] = 0;
disk_mem[19251] = 0;
disk_mem[19252] = 0;
disk_mem[19253] = 0;
disk_mem[19254] = 0;
disk_mem[19255] = 0;
disk_mem[19256] = 0;
disk_mem[19257] = 0;
disk_mem[19258] = 0;
disk_mem[19259] = 0;
disk_mem[19260] = 0;
disk_mem[19261] = 0;
disk_mem[19262] = 0;
disk_mem[19263] = 0;
disk_mem[19264] = 0;
disk_mem[19265] = 0;
disk_mem[19266] = 0;
disk_mem[19267] = 0;
disk_mem[19268] = 0;
disk_mem[19269] = 0;
disk_mem[19270] = 0;
disk_mem[19271] = 0;
disk_mem[19272] = 0;
disk_mem[19273] = 0;
disk_mem[19274] = 0;
disk_mem[19275] = 0;
disk_mem[19276] = 0;
disk_mem[19277] = 0;
disk_mem[19278] = 0;
disk_mem[19279] = 0;
disk_mem[19280] = 0;
disk_mem[19281] = 0;
disk_mem[19282] = 0;
disk_mem[19283] = 0;
disk_mem[19284] = 0;
disk_mem[19285] = 0;
disk_mem[19286] = 0;
disk_mem[19287] = 0;
disk_mem[19288] = 0;
disk_mem[19289] = 0;
disk_mem[19290] = 0;
disk_mem[19291] = 0;
disk_mem[19292] = 0;
disk_mem[19293] = 0;
disk_mem[19294] = 0;
disk_mem[19295] = 0;
disk_mem[19296] = 0;
disk_mem[19297] = 0;
disk_mem[19298] = 0;
disk_mem[19299] = 0;
disk_mem[19300] = 0;
disk_mem[19301] = 0;
disk_mem[19302] = 0;
disk_mem[19303] = 0;
disk_mem[19304] = 0;
disk_mem[19305] = 0;
disk_mem[19306] = 0;
disk_mem[19307] = 0;
disk_mem[19308] = 0;
disk_mem[19309] = 0;
disk_mem[19310] = 0;
disk_mem[19311] = 0;
disk_mem[19312] = 0;
disk_mem[19313] = 0;
disk_mem[19314] = 0;
disk_mem[19315] = 0;
disk_mem[19316] = 0;
disk_mem[19317] = 0;
disk_mem[19318] = 0;
disk_mem[19319] = 0;
disk_mem[19320] = 0;
disk_mem[19321] = 0;
disk_mem[19322] = 0;
disk_mem[19323] = 0;
disk_mem[19324] = 0;
disk_mem[19325] = 0;
disk_mem[19326] = 0;
disk_mem[19327] = 0;
disk_mem[19328] = 0;
disk_mem[19329] = 0;
disk_mem[19330] = 0;
disk_mem[19331] = 0;
disk_mem[19332] = 0;
disk_mem[19333] = 0;
disk_mem[19334] = 0;
disk_mem[19335] = 0;
disk_mem[19336] = 0;
disk_mem[19337] = 0;
disk_mem[19338] = 0;
disk_mem[19339] = 0;
disk_mem[19340] = 0;
disk_mem[19341] = 0;
disk_mem[19342] = 0;
disk_mem[19343] = 0;
disk_mem[19344] = 0;
disk_mem[19345] = 0;
disk_mem[19346] = 0;
disk_mem[19347] = 0;
disk_mem[19348] = 0;
disk_mem[19349] = 0;
disk_mem[19350] = 0;
disk_mem[19351] = 0;
disk_mem[19352] = 0;
disk_mem[19353] = 0;
disk_mem[19354] = 0;
disk_mem[19355] = 0;
disk_mem[19356] = 0;
disk_mem[19357] = 0;
disk_mem[19358] = 0;
disk_mem[19359] = 0;
disk_mem[19360] = 0;
disk_mem[19361] = 0;
disk_mem[19362] = 0;
disk_mem[19363] = 0;
disk_mem[19364] = 0;
disk_mem[19365] = 0;
disk_mem[19366] = 0;
disk_mem[19367] = 0;
disk_mem[19368] = 0;
disk_mem[19369] = 0;
disk_mem[19370] = 0;
disk_mem[19371] = 0;
disk_mem[19372] = 0;
disk_mem[19373] = 0;
disk_mem[19374] = 0;
disk_mem[19375] = 0;
disk_mem[19376] = 0;
disk_mem[19377] = 0;
disk_mem[19378] = 0;
disk_mem[19379] = 0;
disk_mem[19380] = 0;
disk_mem[19381] = 0;
disk_mem[19382] = 0;
disk_mem[19383] = 0;
disk_mem[19384] = 0;
disk_mem[19385] = 0;
disk_mem[19386] = 0;
disk_mem[19387] = 0;
disk_mem[19388] = 0;
disk_mem[19389] = 0;
disk_mem[19390] = 0;
disk_mem[19391] = 0;
disk_mem[19392] = 0;
disk_mem[19393] = 0;
disk_mem[19394] = 0;
disk_mem[19395] = 0;
disk_mem[19396] = 0;
disk_mem[19397] = 0;
disk_mem[19398] = 0;
disk_mem[19399] = 0;
disk_mem[19400] = 0;
disk_mem[19401] = 0;
disk_mem[19402] = 0;
disk_mem[19403] = 0;
disk_mem[19404] = 0;
disk_mem[19405] = 0;
disk_mem[19406] = 0;
disk_mem[19407] = 0;
disk_mem[19408] = 0;
disk_mem[19409] = 0;
disk_mem[19410] = 0;
disk_mem[19411] = 0;
disk_mem[19412] = 0;
disk_mem[19413] = 0;
disk_mem[19414] = 0;
disk_mem[19415] = 0;
disk_mem[19416] = 0;
disk_mem[19417] = 0;
disk_mem[19418] = 0;
disk_mem[19419] = 0;
disk_mem[19420] = 0;
disk_mem[19421] = 0;
disk_mem[19422] = 0;
disk_mem[19423] = 0;
disk_mem[19424] = 0;
disk_mem[19425] = 0;
disk_mem[19426] = 0;
disk_mem[19427] = 0;
disk_mem[19428] = 0;
disk_mem[19429] = 0;
disk_mem[19430] = 0;
disk_mem[19431] = 0;
disk_mem[19432] = 0;
disk_mem[19433] = 0;
disk_mem[19434] = 0;
disk_mem[19435] = 0;
disk_mem[19436] = 0;
disk_mem[19437] = 0;
disk_mem[19438] = 0;
disk_mem[19439] = 0;
disk_mem[19440] = 0;
disk_mem[19441] = 0;
disk_mem[19442] = 0;
disk_mem[19443] = 0;
disk_mem[19444] = 0;
disk_mem[19445] = 0;
disk_mem[19446] = 0;
disk_mem[19447] = 0;
disk_mem[19448] = 0;
disk_mem[19449] = 0;
disk_mem[19450] = 0;
disk_mem[19451] = 0;
disk_mem[19452] = 0;
disk_mem[19453] = 0;
disk_mem[19454] = 0;
disk_mem[19455] = 0;
disk_mem[19456] = 0;
disk_mem[19457] = 0;
disk_mem[19458] = 0;
disk_mem[19459] = 0;
disk_mem[19460] = 0;
disk_mem[19461] = 0;
disk_mem[19462] = 0;
disk_mem[19463] = 0;
disk_mem[19464] = 0;
disk_mem[19465] = 0;
disk_mem[19466] = 0;
disk_mem[19467] = 0;
disk_mem[19468] = 0;
disk_mem[19469] = 0;
disk_mem[19470] = 0;
disk_mem[19471] = 0;
disk_mem[19472] = 0;
disk_mem[19473] = 0;
disk_mem[19474] = 0;
disk_mem[19475] = 0;
disk_mem[19476] = 0;
disk_mem[19477] = 0;
disk_mem[19478] = 0;
disk_mem[19479] = 0;
disk_mem[19480] = 0;
disk_mem[19481] = 0;
disk_mem[19482] = 0;
disk_mem[19483] = 0;
disk_mem[19484] = 0;
disk_mem[19485] = 0;
disk_mem[19486] = 0;
disk_mem[19487] = 0;
disk_mem[19488] = 0;
disk_mem[19489] = 0;
disk_mem[19490] = 0;
disk_mem[19491] = 0;
disk_mem[19492] = 0;
disk_mem[19493] = 0;
disk_mem[19494] = 0;
disk_mem[19495] = 0;
disk_mem[19496] = 0;
disk_mem[19497] = 0;
disk_mem[19498] = 0;
disk_mem[19499] = 0;
disk_mem[19500] = 0;
disk_mem[19501] = 0;
disk_mem[19502] = 0;
disk_mem[19503] = 0;
disk_mem[19504] = 0;
disk_mem[19505] = 0;
disk_mem[19506] = 0;
disk_mem[19507] = 0;
disk_mem[19508] = 0;
disk_mem[19509] = 0;
disk_mem[19510] = 0;
disk_mem[19511] = 0;
disk_mem[19512] = 0;
disk_mem[19513] = 0;
disk_mem[19514] = 0;
disk_mem[19515] = 0;
disk_mem[19516] = 0;
disk_mem[19517] = 0;
disk_mem[19518] = 0;
disk_mem[19519] = 0;
disk_mem[19520] = 0;
disk_mem[19521] = 0;
disk_mem[19522] = 0;
disk_mem[19523] = 0;
disk_mem[19524] = 0;
disk_mem[19525] = 0;
disk_mem[19526] = 0;
disk_mem[19527] = 0;
disk_mem[19528] = 0;
disk_mem[19529] = 0;
disk_mem[19530] = 0;
disk_mem[19531] = 0;
disk_mem[19532] = 0;
disk_mem[19533] = 0;
disk_mem[19534] = 0;
disk_mem[19535] = 0;
disk_mem[19536] = 0;
disk_mem[19537] = 0;
disk_mem[19538] = 0;
disk_mem[19539] = 0;
disk_mem[19540] = 0;
disk_mem[19541] = 0;
disk_mem[19542] = 0;
disk_mem[19543] = 0;
disk_mem[19544] = 0;
disk_mem[19545] = 0;
disk_mem[19546] = 0;
disk_mem[19547] = 0;
disk_mem[19548] = 0;
disk_mem[19549] = 0;
disk_mem[19550] = 0;
disk_mem[19551] = 0;
disk_mem[19552] = 0;
disk_mem[19553] = 0;
disk_mem[19554] = 0;
disk_mem[19555] = 0;
disk_mem[19556] = 0;
disk_mem[19557] = 0;
disk_mem[19558] = 0;
disk_mem[19559] = 0;
disk_mem[19560] = 0;
disk_mem[19561] = 0;
disk_mem[19562] = 0;
disk_mem[19563] = 0;
disk_mem[19564] = 0;
disk_mem[19565] = 0;
disk_mem[19566] = 0;
disk_mem[19567] = 0;
disk_mem[19568] = 0;
disk_mem[19569] = 0;
disk_mem[19570] = 0;
disk_mem[19571] = 0;
disk_mem[19572] = 0;
disk_mem[19573] = 0;
disk_mem[19574] = 0;
disk_mem[19575] = 0;
disk_mem[19576] = 0;
disk_mem[19577] = 0;
disk_mem[19578] = 0;
disk_mem[19579] = 0;
disk_mem[19580] = 0;
disk_mem[19581] = 0;
disk_mem[19582] = 0;
disk_mem[19583] = 0;
disk_mem[19584] = 0;
disk_mem[19585] = 0;
disk_mem[19586] = 0;
disk_mem[19587] = 0;
disk_mem[19588] = 0;
disk_mem[19589] = 0;
disk_mem[19590] = 0;
disk_mem[19591] = 0;
disk_mem[19592] = 0;
disk_mem[19593] = 0;
disk_mem[19594] = 0;
disk_mem[19595] = 0;
disk_mem[19596] = 0;
disk_mem[19597] = 0;
disk_mem[19598] = 0;
disk_mem[19599] = 0;
disk_mem[19600] = 0;
disk_mem[19601] = 0;
disk_mem[19602] = 0;
disk_mem[19603] = 0;
disk_mem[19604] = 0;
disk_mem[19605] = 0;
disk_mem[19606] = 0;
disk_mem[19607] = 0;
disk_mem[19608] = 0;
disk_mem[19609] = 0;
disk_mem[19610] = 0;
disk_mem[19611] = 0;
disk_mem[19612] = 0;
disk_mem[19613] = 0;
disk_mem[19614] = 0;
disk_mem[19615] = 0;
disk_mem[19616] = 0;
disk_mem[19617] = 0;
disk_mem[19618] = 0;
disk_mem[19619] = 0;
disk_mem[19620] = 0;
disk_mem[19621] = 0;
disk_mem[19622] = 0;
disk_mem[19623] = 0;
disk_mem[19624] = 0;
disk_mem[19625] = 0;
disk_mem[19626] = 0;
disk_mem[19627] = 0;
disk_mem[19628] = 0;
disk_mem[19629] = 0;
disk_mem[19630] = 0;
disk_mem[19631] = 0;
disk_mem[19632] = 0;
disk_mem[19633] = 0;
disk_mem[19634] = 0;
disk_mem[19635] = 0;
disk_mem[19636] = 0;
disk_mem[19637] = 0;
disk_mem[19638] = 0;
disk_mem[19639] = 0;
disk_mem[19640] = 0;
disk_mem[19641] = 0;
disk_mem[19642] = 0;
disk_mem[19643] = 0;
disk_mem[19644] = 0;
disk_mem[19645] = 0;
disk_mem[19646] = 0;
disk_mem[19647] = 0;
disk_mem[19648] = 0;
disk_mem[19649] = 0;
disk_mem[19650] = 0;
disk_mem[19651] = 0;
disk_mem[19652] = 0;
disk_mem[19653] = 0;
disk_mem[19654] = 0;
disk_mem[19655] = 0;
disk_mem[19656] = 0;
disk_mem[19657] = 0;
disk_mem[19658] = 0;
disk_mem[19659] = 0;
disk_mem[19660] = 0;
disk_mem[19661] = 0;
disk_mem[19662] = 0;
disk_mem[19663] = 0;
disk_mem[19664] = 0;
disk_mem[19665] = 0;
disk_mem[19666] = 0;
disk_mem[19667] = 0;
disk_mem[19668] = 0;
disk_mem[19669] = 0;
disk_mem[19670] = 0;
disk_mem[19671] = 0;
disk_mem[19672] = 0;
disk_mem[19673] = 0;
disk_mem[19674] = 0;
disk_mem[19675] = 0;
disk_mem[19676] = 0;
disk_mem[19677] = 0;
disk_mem[19678] = 0;
disk_mem[19679] = 0;
disk_mem[19680] = 0;
disk_mem[19681] = 0;
disk_mem[19682] = 0;
disk_mem[19683] = 0;
disk_mem[19684] = 0;
disk_mem[19685] = 0;
disk_mem[19686] = 0;
disk_mem[19687] = 0;
disk_mem[19688] = 0;
disk_mem[19689] = 0;
disk_mem[19690] = 0;
disk_mem[19691] = 0;
disk_mem[19692] = 0;
disk_mem[19693] = 0;
disk_mem[19694] = 0;
disk_mem[19695] = 0;
disk_mem[19696] = 0;
disk_mem[19697] = 0;
disk_mem[19698] = 0;
disk_mem[19699] = 0;
disk_mem[19700] = 0;
disk_mem[19701] = 0;
disk_mem[19702] = 0;
disk_mem[19703] = 0;
disk_mem[19704] = 0;
disk_mem[19705] = 0;
disk_mem[19706] = 0;
disk_mem[19707] = 0;
disk_mem[19708] = 0;
disk_mem[19709] = 0;
disk_mem[19710] = 0;
disk_mem[19711] = 0;
disk_mem[19712] = 0;
disk_mem[19713] = 0;
disk_mem[19714] = 0;
disk_mem[19715] = 0;
disk_mem[19716] = 0;
disk_mem[19717] = 0;
disk_mem[19718] = 0;
disk_mem[19719] = 0;
disk_mem[19720] = 0;
disk_mem[19721] = 0;
disk_mem[19722] = 0;
disk_mem[19723] = 0;
disk_mem[19724] = 0;
disk_mem[19725] = 0;
disk_mem[19726] = 0;
disk_mem[19727] = 0;
disk_mem[19728] = 0;
disk_mem[19729] = 0;
disk_mem[19730] = 0;
disk_mem[19731] = 0;
disk_mem[19732] = 0;
disk_mem[19733] = 0;
disk_mem[19734] = 0;
disk_mem[19735] = 0;
disk_mem[19736] = 0;
disk_mem[19737] = 0;
disk_mem[19738] = 0;
disk_mem[19739] = 0;
disk_mem[19740] = 0;
disk_mem[19741] = 0;
disk_mem[19742] = 0;
disk_mem[19743] = 0;
disk_mem[19744] = 0;
disk_mem[19745] = 0;
disk_mem[19746] = 0;
disk_mem[19747] = 0;
disk_mem[19748] = 0;
disk_mem[19749] = 0;
disk_mem[19750] = 0;
disk_mem[19751] = 0;
disk_mem[19752] = 0;
disk_mem[19753] = 0;
disk_mem[19754] = 0;
disk_mem[19755] = 0;
disk_mem[19756] = 0;
disk_mem[19757] = 0;
disk_mem[19758] = 0;
disk_mem[19759] = 0;
disk_mem[19760] = 0;
disk_mem[19761] = 0;
disk_mem[19762] = 0;
disk_mem[19763] = 0;
disk_mem[19764] = 0;
disk_mem[19765] = 0;
disk_mem[19766] = 0;
disk_mem[19767] = 0;
disk_mem[19768] = 0;
disk_mem[19769] = 0;
disk_mem[19770] = 0;
disk_mem[19771] = 0;
disk_mem[19772] = 0;
disk_mem[19773] = 0;
disk_mem[19774] = 0;
disk_mem[19775] = 0;
disk_mem[19776] = 0;
disk_mem[19777] = 0;
disk_mem[19778] = 0;
disk_mem[19779] = 0;
disk_mem[19780] = 0;
disk_mem[19781] = 0;
disk_mem[19782] = 0;
disk_mem[19783] = 0;
disk_mem[19784] = 0;
disk_mem[19785] = 0;
disk_mem[19786] = 0;
disk_mem[19787] = 0;
disk_mem[19788] = 0;
disk_mem[19789] = 0;
disk_mem[19790] = 0;
disk_mem[19791] = 0;
disk_mem[19792] = 0;
disk_mem[19793] = 0;
disk_mem[19794] = 0;
disk_mem[19795] = 0;
disk_mem[19796] = 0;
disk_mem[19797] = 0;
disk_mem[19798] = 0;
disk_mem[19799] = 0;
disk_mem[19800] = 0;
disk_mem[19801] = 0;
disk_mem[19802] = 0;
disk_mem[19803] = 0;
disk_mem[19804] = 0;
disk_mem[19805] = 0;
disk_mem[19806] = 0;
disk_mem[19807] = 0;
disk_mem[19808] = 0;
disk_mem[19809] = 0;
disk_mem[19810] = 0;
disk_mem[19811] = 0;
disk_mem[19812] = 0;
disk_mem[19813] = 0;
disk_mem[19814] = 0;
disk_mem[19815] = 0;
disk_mem[19816] = 0;
disk_mem[19817] = 0;
disk_mem[19818] = 0;
disk_mem[19819] = 0;
disk_mem[19820] = 0;
disk_mem[19821] = 0;
disk_mem[19822] = 0;
disk_mem[19823] = 0;
disk_mem[19824] = 0;
disk_mem[19825] = 0;
disk_mem[19826] = 0;
disk_mem[19827] = 0;
disk_mem[19828] = 0;
disk_mem[19829] = 0;
disk_mem[19830] = 0;
disk_mem[19831] = 0;
disk_mem[19832] = 0;
disk_mem[19833] = 0;
disk_mem[19834] = 0;
disk_mem[19835] = 0;
disk_mem[19836] = 0;
disk_mem[19837] = 0;
disk_mem[19838] = 0;
disk_mem[19839] = 0;
disk_mem[19840] = 0;
disk_mem[19841] = 0;
disk_mem[19842] = 0;
disk_mem[19843] = 0;
disk_mem[19844] = 0;
disk_mem[19845] = 0;
disk_mem[19846] = 0;
disk_mem[19847] = 0;
disk_mem[19848] = 0;
disk_mem[19849] = 0;
disk_mem[19850] = 0;
disk_mem[19851] = 0;
disk_mem[19852] = 0;
disk_mem[19853] = 0;
disk_mem[19854] = 0;
disk_mem[19855] = 0;
disk_mem[19856] = 0;
disk_mem[19857] = 0;
disk_mem[19858] = 0;
disk_mem[19859] = 0;
disk_mem[19860] = 0;
disk_mem[19861] = 0;
disk_mem[19862] = 0;
disk_mem[19863] = 0;
disk_mem[19864] = 0;
disk_mem[19865] = 0;
disk_mem[19866] = 0;
disk_mem[19867] = 0;
disk_mem[19868] = 0;
disk_mem[19869] = 0;
disk_mem[19870] = 0;
disk_mem[19871] = 0;
disk_mem[19872] = 0;
disk_mem[19873] = 0;
disk_mem[19874] = 0;
disk_mem[19875] = 0;
disk_mem[19876] = 0;
disk_mem[19877] = 0;
disk_mem[19878] = 0;
disk_mem[19879] = 0;
disk_mem[19880] = 0;
disk_mem[19881] = 0;
disk_mem[19882] = 0;
disk_mem[19883] = 0;
disk_mem[19884] = 0;
disk_mem[19885] = 0;
disk_mem[19886] = 0;
disk_mem[19887] = 0;
disk_mem[19888] = 0;
disk_mem[19889] = 0;
disk_mem[19890] = 0;
disk_mem[19891] = 0;
disk_mem[19892] = 0;
disk_mem[19893] = 0;
disk_mem[19894] = 0;
disk_mem[19895] = 0;
disk_mem[19896] = 0;
disk_mem[19897] = 0;
disk_mem[19898] = 0;
disk_mem[19899] = 0;
disk_mem[19900] = 0;
disk_mem[19901] = 0;
disk_mem[19902] = 0;
disk_mem[19903] = 0;
disk_mem[19904] = 0;
disk_mem[19905] = 0;
disk_mem[19906] = 0;
disk_mem[19907] = 0;
disk_mem[19908] = 0;
disk_mem[19909] = 0;
disk_mem[19910] = 0;
disk_mem[19911] = 0;
disk_mem[19912] = 0;
disk_mem[19913] = 0;
disk_mem[19914] = 0;
disk_mem[19915] = 0;
disk_mem[19916] = 0;
disk_mem[19917] = 0;
disk_mem[19918] = 0;
disk_mem[19919] = 0;
disk_mem[19920] = 0;
disk_mem[19921] = 0;
disk_mem[19922] = 0;
disk_mem[19923] = 0;
disk_mem[19924] = 0;
disk_mem[19925] = 0;
disk_mem[19926] = 0;
disk_mem[19927] = 0;
disk_mem[19928] = 0;
disk_mem[19929] = 0;
disk_mem[19930] = 0;
disk_mem[19931] = 0;
disk_mem[19932] = 0;
disk_mem[19933] = 0;
disk_mem[19934] = 0;
disk_mem[19935] = 0;
disk_mem[19936] = 0;
disk_mem[19937] = 0;
disk_mem[19938] = 0;
disk_mem[19939] = 0;
disk_mem[19940] = 0;
disk_mem[19941] = 0;
disk_mem[19942] = 0;
disk_mem[19943] = 0;
disk_mem[19944] = 0;
disk_mem[19945] = 0;
disk_mem[19946] = 0;
disk_mem[19947] = 0;
disk_mem[19948] = 0;
disk_mem[19949] = 0;
disk_mem[19950] = 0;
disk_mem[19951] = 0;
disk_mem[19952] = 0;
disk_mem[19953] = 0;
disk_mem[19954] = 0;
disk_mem[19955] = 0;
disk_mem[19956] = 0;
disk_mem[19957] = 0;
disk_mem[19958] = 0;
disk_mem[19959] = 0;
disk_mem[19960] = 0;
disk_mem[19961] = 0;
disk_mem[19962] = 0;
disk_mem[19963] = 0;
disk_mem[19964] = 0;
disk_mem[19965] = 0;
disk_mem[19966] = 0;
disk_mem[19967] = 0;
disk_mem[19968] = 0;
disk_mem[19969] = 0;
disk_mem[19970] = 0;
disk_mem[19971] = 0;
disk_mem[19972] = 0;
disk_mem[19973] = 0;
disk_mem[19974] = 0;
disk_mem[19975] = 0;
disk_mem[19976] = 0;
disk_mem[19977] = 0;
disk_mem[19978] = 0;
disk_mem[19979] = 0;
disk_mem[19980] = 0;
disk_mem[19981] = 0;
disk_mem[19982] = 0;
disk_mem[19983] = 0;
disk_mem[19984] = 0;
disk_mem[19985] = 0;
disk_mem[19986] = 0;
disk_mem[19987] = 0;
disk_mem[19988] = 0;
disk_mem[19989] = 0;
disk_mem[19990] = 0;
disk_mem[19991] = 0;
disk_mem[19992] = 0;
disk_mem[19993] = 0;
disk_mem[19994] = 0;
disk_mem[19995] = 0;
disk_mem[19996] = 0;
disk_mem[19997] = 0;
disk_mem[19998] = 0;
disk_mem[19999] = 0;
disk_mem[20000] = 0;
disk_mem[20001] = 0;
disk_mem[20002] = 0;
disk_mem[20003] = 0;
disk_mem[20004] = 0;
disk_mem[20005] = 0;
disk_mem[20006] = 0;
disk_mem[20007] = 0;
disk_mem[20008] = 0;
disk_mem[20009] = 0;
disk_mem[20010] = 0;
disk_mem[20011] = 0;
disk_mem[20012] = 0;
disk_mem[20013] = 0;
disk_mem[20014] = 0;
disk_mem[20015] = 0;
disk_mem[20016] = 0;
disk_mem[20017] = 0;
disk_mem[20018] = 0;
disk_mem[20019] = 0;
disk_mem[20020] = 0;
disk_mem[20021] = 0;
disk_mem[20022] = 0;
disk_mem[20023] = 0;
disk_mem[20024] = 0;
disk_mem[20025] = 0;
disk_mem[20026] = 0;
disk_mem[20027] = 0;
disk_mem[20028] = 0;
disk_mem[20029] = 0;
disk_mem[20030] = 0;
disk_mem[20031] = 0;
disk_mem[20032] = 0;
disk_mem[20033] = 0;
disk_mem[20034] = 0;
disk_mem[20035] = 0;
disk_mem[20036] = 0;
disk_mem[20037] = 0;
disk_mem[20038] = 0;
disk_mem[20039] = 0;
disk_mem[20040] = 0;
disk_mem[20041] = 0;
disk_mem[20042] = 0;
disk_mem[20043] = 0;
disk_mem[20044] = 0;
disk_mem[20045] = 0;
disk_mem[20046] = 0;
disk_mem[20047] = 0;
disk_mem[20048] = 0;
disk_mem[20049] = 0;
disk_mem[20050] = 0;
disk_mem[20051] = 0;
disk_mem[20052] = 0;
disk_mem[20053] = 0;
disk_mem[20054] = 0;
disk_mem[20055] = 0;
disk_mem[20056] = 0;
disk_mem[20057] = 0;
disk_mem[20058] = 0;
disk_mem[20059] = 0;
disk_mem[20060] = 0;
disk_mem[20061] = 0;
disk_mem[20062] = 0;
disk_mem[20063] = 0;
disk_mem[20064] = 0;
disk_mem[20065] = 0;
disk_mem[20066] = 0;
disk_mem[20067] = 0;
disk_mem[20068] = 0;
disk_mem[20069] = 0;
disk_mem[20070] = 0;
disk_mem[20071] = 0;
disk_mem[20072] = 0;
disk_mem[20073] = 0;
disk_mem[20074] = 0;
disk_mem[20075] = 0;
disk_mem[20076] = 0;
disk_mem[20077] = 0;
disk_mem[20078] = 0;
disk_mem[20079] = 0;
disk_mem[20080] = 0;
disk_mem[20081] = 0;
disk_mem[20082] = 0;
disk_mem[20083] = 0;
disk_mem[20084] = 0;
disk_mem[20085] = 0;
disk_mem[20086] = 0;
disk_mem[20087] = 0;
disk_mem[20088] = 0;
disk_mem[20089] = 0;
disk_mem[20090] = 0;
disk_mem[20091] = 0;
disk_mem[20092] = 0;
disk_mem[20093] = 0;
disk_mem[20094] = 0;
disk_mem[20095] = 0;
disk_mem[20096] = 0;
disk_mem[20097] = 0;
disk_mem[20098] = 0;
disk_mem[20099] = 0;
disk_mem[20100] = 0;
disk_mem[20101] = 0;
disk_mem[20102] = 0;
disk_mem[20103] = 0;
disk_mem[20104] = 0;
disk_mem[20105] = 0;
disk_mem[20106] = 0;
disk_mem[20107] = 0;
disk_mem[20108] = 0;
disk_mem[20109] = 0;
disk_mem[20110] = 0;
disk_mem[20111] = 0;
disk_mem[20112] = 0;
disk_mem[20113] = 0;
disk_mem[20114] = 0;
disk_mem[20115] = 0;
disk_mem[20116] = 0;
disk_mem[20117] = 0;
disk_mem[20118] = 0;
disk_mem[20119] = 0;
disk_mem[20120] = 0;
disk_mem[20121] = 0;
disk_mem[20122] = 0;
disk_mem[20123] = 0;
disk_mem[20124] = 0;
disk_mem[20125] = 0;
disk_mem[20126] = 0;
disk_mem[20127] = 0;
disk_mem[20128] = 0;
disk_mem[20129] = 0;
disk_mem[20130] = 0;
disk_mem[20131] = 0;
disk_mem[20132] = 0;
disk_mem[20133] = 0;
disk_mem[20134] = 0;
disk_mem[20135] = 0;
disk_mem[20136] = 0;
disk_mem[20137] = 0;
disk_mem[20138] = 0;
disk_mem[20139] = 0;
disk_mem[20140] = 0;
disk_mem[20141] = 0;
disk_mem[20142] = 0;
disk_mem[20143] = 0;
disk_mem[20144] = 0;
disk_mem[20145] = 0;
disk_mem[20146] = 0;
disk_mem[20147] = 0;
disk_mem[20148] = 0;
disk_mem[20149] = 0;
disk_mem[20150] = 0;
disk_mem[20151] = 0;
disk_mem[20152] = 0;
disk_mem[20153] = 0;
disk_mem[20154] = 0;
disk_mem[20155] = 0;
disk_mem[20156] = 0;
disk_mem[20157] = 0;
disk_mem[20158] = 0;
disk_mem[20159] = 0;
disk_mem[20160] = 0;
disk_mem[20161] = 0;
disk_mem[20162] = 0;
disk_mem[20163] = 0;
disk_mem[20164] = 0;
disk_mem[20165] = 0;
disk_mem[20166] = 0;
disk_mem[20167] = 0;
disk_mem[20168] = 0;
disk_mem[20169] = 0;
disk_mem[20170] = 0;
disk_mem[20171] = 0;
disk_mem[20172] = 0;
disk_mem[20173] = 0;
disk_mem[20174] = 0;
disk_mem[20175] = 0;
disk_mem[20176] = 0;
disk_mem[20177] = 0;
disk_mem[20178] = 0;
disk_mem[20179] = 0;
disk_mem[20180] = 0;
disk_mem[20181] = 0;
disk_mem[20182] = 0;
disk_mem[20183] = 0;
disk_mem[20184] = 0;
disk_mem[20185] = 0;
disk_mem[20186] = 0;
disk_mem[20187] = 0;
disk_mem[20188] = 0;
disk_mem[20189] = 0;
disk_mem[20190] = 0;
disk_mem[20191] = 0;
disk_mem[20192] = 0;
disk_mem[20193] = 0;
disk_mem[20194] = 0;
disk_mem[20195] = 0;
disk_mem[20196] = 0;
disk_mem[20197] = 0;
disk_mem[20198] = 0;
disk_mem[20199] = 0;
disk_mem[20200] = 0;
disk_mem[20201] = 0;
disk_mem[20202] = 0;
disk_mem[20203] = 0;
disk_mem[20204] = 0;
disk_mem[20205] = 0;
disk_mem[20206] = 0;
disk_mem[20207] = 0;
disk_mem[20208] = 0;
disk_mem[20209] = 0;
disk_mem[20210] = 0;
disk_mem[20211] = 0;
disk_mem[20212] = 0;
disk_mem[20213] = 0;
disk_mem[20214] = 0;
disk_mem[20215] = 0;
disk_mem[20216] = 0;
disk_mem[20217] = 0;
disk_mem[20218] = 0;
disk_mem[20219] = 0;
disk_mem[20220] = 0;
disk_mem[20221] = 0;
disk_mem[20222] = 0;
disk_mem[20223] = 0;
disk_mem[20224] = 0;
disk_mem[20225] = 0;
disk_mem[20226] = 0;
disk_mem[20227] = 0;
disk_mem[20228] = 0;
disk_mem[20229] = 0;
disk_mem[20230] = 0;
disk_mem[20231] = 0;
disk_mem[20232] = 0;
disk_mem[20233] = 0;
disk_mem[20234] = 0;
disk_mem[20235] = 0;
disk_mem[20236] = 0;
disk_mem[20237] = 0;
disk_mem[20238] = 0;
disk_mem[20239] = 0;
disk_mem[20240] = 0;
disk_mem[20241] = 0;
disk_mem[20242] = 0;
disk_mem[20243] = 0;
disk_mem[20244] = 0;
disk_mem[20245] = 0;
disk_mem[20246] = 0;
disk_mem[20247] = 0;
disk_mem[20248] = 0;
disk_mem[20249] = 0;
disk_mem[20250] = 0;
disk_mem[20251] = 0;
disk_mem[20252] = 0;
disk_mem[20253] = 0;
disk_mem[20254] = 0;
disk_mem[20255] = 0;
disk_mem[20256] = 0;
disk_mem[20257] = 0;
disk_mem[20258] = 0;
disk_mem[20259] = 0;
disk_mem[20260] = 0;
disk_mem[20261] = 0;
disk_mem[20262] = 0;
disk_mem[20263] = 0;
disk_mem[20264] = 0;
disk_mem[20265] = 0;
disk_mem[20266] = 0;
disk_mem[20267] = 0;
disk_mem[20268] = 0;
disk_mem[20269] = 0;
disk_mem[20270] = 0;
disk_mem[20271] = 0;
disk_mem[20272] = 0;
disk_mem[20273] = 0;
disk_mem[20274] = 0;
disk_mem[20275] = 0;
disk_mem[20276] = 0;
disk_mem[20277] = 0;
disk_mem[20278] = 0;
disk_mem[20279] = 0;
disk_mem[20280] = 0;
disk_mem[20281] = 0;
disk_mem[20282] = 0;
disk_mem[20283] = 0;
disk_mem[20284] = 0;
disk_mem[20285] = 0;
disk_mem[20286] = 0;
disk_mem[20287] = 0;
disk_mem[20288] = 0;
disk_mem[20289] = 0;
disk_mem[20290] = 0;
disk_mem[20291] = 0;
disk_mem[20292] = 0;
disk_mem[20293] = 0;
disk_mem[20294] = 0;
disk_mem[20295] = 0;
disk_mem[20296] = 0;
disk_mem[20297] = 0;
disk_mem[20298] = 0;
disk_mem[20299] = 0;
disk_mem[20300] = 0;
disk_mem[20301] = 0;
disk_mem[20302] = 0;
disk_mem[20303] = 0;
disk_mem[20304] = 0;
disk_mem[20305] = 0;
disk_mem[20306] = 0;
disk_mem[20307] = 0;
disk_mem[20308] = 0;
disk_mem[20309] = 0;
disk_mem[20310] = 0;
disk_mem[20311] = 0;
disk_mem[20312] = 0;
disk_mem[20313] = 0;
disk_mem[20314] = 0;
disk_mem[20315] = 0;
disk_mem[20316] = 0;
disk_mem[20317] = 0;
disk_mem[20318] = 0;
disk_mem[20319] = 0;
disk_mem[20320] = 0;
disk_mem[20321] = 0;
disk_mem[20322] = 0;
disk_mem[20323] = 0;
disk_mem[20324] = 0;
disk_mem[20325] = 0;
disk_mem[20326] = 0;
disk_mem[20327] = 0;
disk_mem[20328] = 0;
disk_mem[20329] = 0;
disk_mem[20330] = 0;
disk_mem[20331] = 0;
disk_mem[20332] = 0;
disk_mem[20333] = 0;
disk_mem[20334] = 0;
disk_mem[20335] = 0;
disk_mem[20336] = 0;
disk_mem[20337] = 0;
disk_mem[20338] = 0;
disk_mem[20339] = 0;
disk_mem[20340] = 0;
disk_mem[20341] = 0;
disk_mem[20342] = 0;
disk_mem[20343] = 0;
disk_mem[20344] = 0;
disk_mem[20345] = 0;
disk_mem[20346] = 0;
disk_mem[20347] = 0;
disk_mem[20348] = 0;
disk_mem[20349] = 0;
disk_mem[20350] = 0;
disk_mem[20351] = 0;
disk_mem[20352] = 0;
disk_mem[20353] = 0;
disk_mem[20354] = 0;
disk_mem[20355] = 0;
disk_mem[20356] = 0;
disk_mem[20357] = 0;
disk_mem[20358] = 0;
disk_mem[20359] = 0;
disk_mem[20360] = 0;
disk_mem[20361] = 0;
disk_mem[20362] = 0;
disk_mem[20363] = 0;
disk_mem[20364] = 0;
disk_mem[20365] = 0;
disk_mem[20366] = 0;
disk_mem[20367] = 0;
disk_mem[20368] = 0;
disk_mem[20369] = 0;
disk_mem[20370] = 0;
disk_mem[20371] = 0;
disk_mem[20372] = 0;
disk_mem[20373] = 0;
disk_mem[20374] = 0;
disk_mem[20375] = 0;
disk_mem[20376] = 0;
disk_mem[20377] = 0;
disk_mem[20378] = 0;
disk_mem[20379] = 0;
disk_mem[20380] = 0;
disk_mem[20381] = 0;
disk_mem[20382] = 0;
disk_mem[20383] = 0;
disk_mem[20384] = 0;
disk_mem[20385] = 0;
disk_mem[20386] = 0;
disk_mem[20387] = 0;
disk_mem[20388] = 0;
disk_mem[20389] = 0;
disk_mem[20390] = 0;
disk_mem[20391] = 0;
disk_mem[20392] = 0;
disk_mem[20393] = 0;
disk_mem[20394] = 0;
disk_mem[20395] = 0;
disk_mem[20396] = 0;
disk_mem[20397] = 0;
disk_mem[20398] = 0;
disk_mem[20399] = 0;
disk_mem[20400] = 0;
disk_mem[20401] = 0;
disk_mem[20402] = 0;
disk_mem[20403] = 0;
disk_mem[20404] = 0;
disk_mem[20405] = 0;
disk_mem[20406] = 0;
disk_mem[20407] = 0;
disk_mem[20408] = 0;
disk_mem[20409] = 0;
disk_mem[20410] = 0;
disk_mem[20411] = 0;
disk_mem[20412] = 0;
disk_mem[20413] = 0;
disk_mem[20414] = 0;
disk_mem[20415] = 0;
disk_mem[20416] = 0;
disk_mem[20417] = 0;
disk_mem[20418] = 0;
disk_mem[20419] = 0;
disk_mem[20420] = 0;
disk_mem[20421] = 0;
disk_mem[20422] = 0;
disk_mem[20423] = 0;
disk_mem[20424] = 0;
disk_mem[20425] = 0;
disk_mem[20426] = 0;
disk_mem[20427] = 0;
disk_mem[20428] = 0;
disk_mem[20429] = 0;
disk_mem[20430] = 0;
disk_mem[20431] = 0;
disk_mem[20432] = 0;
disk_mem[20433] = 0;
disk_mem[20434] = 0;
disk_mem[20435] = 0;
disk_mem[20436] = 0;
disk_mem[20437] = 0;
disk_mem[20438] = 0;
disk_mem[20439] = 0;
disk_mem[20440] = 0;
disk_mem[20441] = 0;
disk_mem[20442] = 0;
disk_mem[20443] = 0;
disk_mem[20444] = 0;
disk_mem[20445] = 0;
disk_mem[20446] = 0;
disk_mem[20447] = 0;
disk_mem[20448] = 0;
disk_mem[20449] = 0;
disk_mem[20450] = 0;
disk_mem[20451] = 0;
disk_mem[20452] = 0;
disk_mem[20453] = 0;
disk_mem[20454] = 0;
disk_mem[20455] = 0;
disk_mem[20456] = 0;
disk_mem[20457] = 0;
disk_mem[20458] = 0;
disk_mem[20459] = 0;
disk_mem[20460] = 0;
disk_mem[20461] = 0;
disk_mem[20462] = 0;
disk_mem[20463] = 0;
disk_mem[20464] = 0;
disk_mem[20465] = 0;
disk_mem[20466] = 0;
disk_mem[20467] = 0;
disk_mem[20468] = 0;
disk_mem[20469] = 0;
disk_mem[20470] = 0;
disk_mem[20471] = 0;
disk_mem[20472] = 0;
disk_mem[20473] = 0;
disk_mem[20474] = 0;
disk_mem[20475] = 0;
disk_mem[20476] = 0;
disk_mem[20477] = 0;
disk_mem[20478] = 0;
disk_mem[20479] = 0;
disk_mem[20480] = 0;
disk_mem[20481] = 0;
disk_mem[20482] = 0;
disk_mem[20483] = 0;
disk_mem[20484] = 0;
disk_mem[20485] = 0;
disk_mem[20486] = 0;
disk_mem[20487] = 0;
disk_mem[20488] = 0;
disk_mem[20489] = 0;
disk_mem[20490] = 0;
disk_mem[20491] = 0;
disk_mem[20492] = 0;
disk_mem[20493] = 0;
disk_mem[20494] = 0;
disk_mem[20495] = 0;
disk_mem[20496] = 0;
disk_mem[20497] = 0;
disk_mem[20498] = 0;
disk_mem[20499] = 0;
disk_mem[20500] = 0;
disk_mem[20501] = 0;
disk_mem[20502] = 0;
disk_mem[20503] = 0;
disk_mem[20504] = 0;
disk_mem[20505] = 0;
disk_mem[20506] = 0;
disk_mem[20507] = 0;
disk_mem[20508] = 0;
disk_mem[20509] = 0;
disk_mem[20510] = 0;
disk_mem[20511] = 0;
disk_mem[20512] = 0;
disk_mem[20513] = 0;
disk_mem[20514] = 0;
disk_mem[20515] = 0;
disk_mem[20516] = 0;
disk_mem[20517] = 0;
disk_mem[20518] = 0;
disk_mem[20519] = 0;
disk_mem[20520] = 0;
disk_mem[20521] = 0;
disk_mem[20522] = 0;
disk_mem[20523] = 0;
disk_mem[20524] = 0;
disk_mem[20525] = 0;
disk_mem[20526] = 0;
disk_mem[20527] = 0;
disk_mem[20528] = 0;
disk_mem[20529] = 0;
disk_mem[20530] = 0;
disk_mem[20531] = 0;
disk_mem[20532] = 0;
disk_mem[20533] = 0;
disk_mem[20534] = 0;
disk_mem[20535] = 0;
disk_mem[20536] = 0;
disk_mem[20537] = 0;
disk_mem[20538] = 0;
disk_mem[20539] = 0;
disk_mem[20540] = 0;
disk_mem[20541] = 0;
disk_mem[20542] = 0;
disk_mem[20543] = 0;
disk_mem[20544] = 0;
disk_mem[20545] = 0;
disk_mem[20546] = 0;
disk_mem[20547] = 0;
disk_mem[20548] = 0;
disk_mem[20549] = 0;
disk_mem[20550] = 0;
disk_mem[20551] = 0;
disk_mem[20552] = 0;
disk_mem[20553] = 0;
disk_mem[20554] = 0;
disk_mem[20555] = 0;
disk_mem[20556] = 0;
disk_mem[20557] = 0;
disk_mem[20558] = 0;
disk_mem[20559] = 0;
disk_mem[20560] = 0;
disk_mem[20561] = 0;
disk_mem[20562] = 0;
disk_mem[20563] = 0;
disk_mem[20564] = 0;
disk_mem[20565] = 0;
disk_mem[20566] = 0;
disk_mem[20567] = 0;
disk_mem[20568] = 0;
disk_mem[20569] = 0;
disk_mem[20570] = 0;
disk_mem[20571] = 0;
disk_mem[20572] = 0;
disk_mem[20573] = 0;
disk_mem[20574] = 0;
disk_mem[20575] = 0;
disk_mem[20576] = 0;
disk_mem[20577] = 0;
disk_mem[20578] = 0;
disk_mem[20579] = 0;
disk_mem[20580] = 0;
disk_mem[20581] = 0;
disk_mem[20582] = 0;
disk_mem[20583] = 0;
disk_mem[20584] = 0;
disk_mem[20585] = 0;
disk_mem[20586] = 0;
disk_mem[20587] = 0;
disk_mem[20588] = 0;
disk_mem[20589] = 0;
disk_mem[20590] = 0;
disk_mem[20591] = 0;
disk_mem[20592] = 0;
disk_mem[20593] = 0;
disk_mem[20594] = 0;
disk_mem[20595] = 0;
disk_mem[20596] = 0;
disk_mem[20597] = 0;
disk_mem[20598] = 0;
disk_mem[20599] = 0;
disk_mem[20600] = 0;
disk_mem[20601] = 0;
disk_mem[20602] = 0;
disk_mem[20603] = 0;
disk_mem[20604] = 0;
disk_mem[20605] = 0;
disk_mem[20606] = 0;
disk_mem[20607] = 0;
disk_mem[20608] = 0;
disk_mem[20609] = 0;
disk_mem[20610] = 0;
disk_mem[20611] = 0;
disk_mem[20612] = 0;
disk_mem[20613] = 0;
disk_mem[20614] = 0;
disk_mem[20615] = 0;
disk_mem[20616] = 0;
disk_mem[20617] = 0;
disk_mem[20618] = 0;
disk_mem[20619] = 0;
disk_mem[20620] = 0;
disk_mem[20621] = 0;
disk_mem[20622] = 0;
disk_mem[20623] = 0;
disk_mem[20624] = 0;
disk_mem[20625] = 0;
disk_mem[20626] = 0;
disk_mem[20627] = 0;
disk_mem[20628] = 0;
disk_mem[20629] = 0;
disk_mem[20630] = 0;
disk_mem[20631] = 0;
disk_mem[20632] = 0;
disk_mem[20633] = 0;
disk_mem[20634] = 0;
disk_mem[20635] = 0;
disk_mem[20636] = 0;
disk_mem[20637] = 0;
disk_mem[20638] = 0;
disk_mem[20639] = 0;
disk_mem[20640] = 0;
disk_mem[20641] = 0;
disk_mem[20642] = 0;
disk_mem[20643] = 0;
disk_mem[20644] = 0;
disk_mem[20645] = 0;
disk_mem[20646] = 0;
disk_mem[20647] = 0;
disk_mem[20648] = 0;
disk_mem[20649] = 0;
disk_mem[20650] = 0;
disk_mem[20651] = 0;
disk_mem[20652] = 0;
disk_mem[20653] = 0;
disk_mem[20654] = 0;
disk_mem[20655] = 0;
disk_mem[20656] = 0;
disk_mem[20657] = 0;
disk_mem[20658] = 0;
disk_mem[20659] = 0;
disk_mem[20660] = 0;
disk_mem[20661] = 0;
disk_mem[20662] = 0;
disk_mem[20663] = 0;
disk_mem[20664] = 0;
disk_mem[20665] = 0;
disk_mem[20666] = 0;
disk_mem[20667] = 0;
disk_mem[20668] = 0;
disk_mem[20669] = 0;
disk_mem[20670] = 0;
disk_mem[20671] = 0;
disk_mem[20672] = 0;
disk_mem[20673] = 0;
disk_mem[20674] = 0;
disk_mem[20675] = 0;
disk_mem[20676] = 0;
disk_mem[20677] = 0;
disk_mem[20678] = 0;
disk_mem[20679] = 0;
disk_mem[20680] = 0;
disk_mem[20681] = 0;
disk_mem[20682] = 0;
disk_mem[20683] = 0;
disk_mem[20684] = 0;
disk_mem[20685] = 0;
disk_mem[20686] = 0;
disk_mem[20687] = 0;
disk_mem[20688] = 0;
disk_mem[20689] = 0;
disk_mem[20690] = 0;
disk_mem[20691] = 0;
disk_mem[20692] = 0;
disk_mem[20693] = 0;
disk_mem[20694] = 0;
disk_mem[20695] = 0;
disk_mem[20696] = 0;
disk_mem[20697] = 0;
disk_mem[20698] = 0;
disk_mem[20699] = 0;
disk_mem[20700] = 0;
disk_mem[20701] = 0;
disk_mem[20702] = 0;
disk_mem[20703] = 0;
disk_mem[20704] = 0;
disk_mem[20705] = 0;
disk_mem[20706] = 0;
disk_mem[20707] = 0;
disk_mem[20708] = 0;
disk_mem[20709] = 0;
disk_mem[20710] = 0;
disk_mem[20711] = 0;
disk_mem[20712] = 0;
disk_mem[20713] = 0;
disk_mem[20714] = 0;
disk_mem[20715] = 0;
disk_mem[20716] = 0;
disk_mem[20717] = 0;
disk_mem[20718] = 0;
disk_mem[20719] = 0;
disk_mem[20720] = 0;
disk_mem[20721] = 0;
disk_mem[20722] = 0;
disk_mem[20723] = 0;
disk_mem[20724] = 0;
disk_mem[20725] = 0;
disk_mem[20726] = 0;
disk_mem[20727] = 0;
disk_mem[20728] = 0;
disk_mem[20729] = 0;
disk_mem[20730] = 0;
disk_mem[20731] = 0;
disk_mem[20732] = 0;
disk_mem[20733] = 0;
disk_mem[20734] = 0;
disk_mem[20735] = 0;
disk_mem[20736] = 0;
disk_mem[20737] = 0;
disk_mem[20738] = 0;
disk_mem[20739] = 0;
disk_mem[20740] = 0;
disk_mem[20741] = 0;
disk_mem[20742] = 0;
disk_mem[20743] = 0;
disk_mem[20744] = 0;
disk_mem[20745] = 0;
disk_mem[20746] = 0;
disk_mem[20747] = 0;
disk_mem[20748] = 0;
disk_mem[20749] = 0;
disk_mem[20750] = 0;
disk_mem[20751] = 0;
disk_mem[20752] = 0;
disk_mem[20753] = 0;
disk_mem[20754] = 0;
disk_mem[20755] = 0;
disk_mem[20756] = 0;
disk_mem[20757] = 0;
disk_mem[20758] = 0;
disk_mem[20759] = 0;
disk_mem[20760] = 0;
disk_mem[20761] = 0;
disk_mem[20762] = 0;
disk_mem[20763] = 0;
disk_mem[20764] = 0;
disk_mem[20765] = 0;
disk_mem[20766] = 0;
disk_mem[20767] = 0;
disk_mem[20768] = 0;
disk_mem[20769] = 0;
disk_mem[20770] = 0;
disk_mem[20771] = 0;
disk_mem[20772] = 0;
disk_mem[20773] = 0;
disk_mem[20774] = 0;
disk_mem[20775] = 0;
disk_mem[20776] = 0;
disk_mem[20777] = 0;
disk_mem[20778] = 0;
disk_mem[20779] = 0;
disk_mem[20780] = 0;
disk_mem[20781] = 0;
disk_mem[20782] = 0;
disk_mem[20783] = 0;
disk_mem[20784] = 0;
disk_mem[20785] = 0;
disk_mem[20786] = 0;
disk_mem[20787] = 0;
disk_mem[20788] = 0;
disk_mem[20789] = 0;
disk_mem[20790] = 0;
disk_mem[20791] = 0;
disk_mem[20792] = 0;
disk_mem[20793] = 0;
disk_mem[20794] = 0;
disk_mem[20795] = 0;
disk_mem[20796] = 0;
disk_mem[20797] = 0;
disk_mem[20798] = 0;
disk_mem[20799] = 0;
disk_mem[20800] = 0;
disk_mem[20801] = 0;
disk_mem[20802] = 0;
disk_mem[20803] = 0;
disk_mem[20804] = 0;
disk_mem[20805] = 0;
disk_mem[20806] = 0;
disk_mem[20807] = 0;
disk_mem[20808] = 0;
disk_mem[20809] = 0;
disk_mem[20810] = 0;
disk_mem[20811] = 0;
disk_mem[20812] = 0;
disk_mem[20813] = 0;
disk_mem[20814] = 0;
disk_mem[20815] = 0;
disk_mem[20816] = 0;
disk_mem[20817] = 0;
disk_mem[20818] = 0;
disk_mem[20819] = 0;
disk_mem[20820] = 0;
disk_mem[20821] = 0;
disk_mem[20822] = 0;
disk_mem[20823] = 0;
disk_mem[20824] = 0;
disk_mem[20825] = 0;
disk_mem[20826] = 0;
disk_mem[20827] = 0;
disk_mem[20828] = 0;
disk_mem[20829] = 0;
disk_mem[20830] = 0;
disk_mem[20831] = 0;
disk_mem[20832] = 0;
disk_mem[20833] = 0;
disk_mem[20834] = 0;
disk_mem[20835] = 0;
disk_mem[20836] = 0;
disk_mem[20837] = 0;
disk_mem[20838] = 0;
disk_mem[20839] = 0;
disk_mem[20840] = 0;
disk_mem[20841] = 0;
disk_mem[20842] = 0;
disk_mem[20843] = 0;
disk_mem[20844] = 0;
disk_mem[20845] = 0;
disk_mem[20846] = 0;
disk_mem[20847] = 0;
disk_mem[20848] = 0;
disk_mem[20849] = 0;
disk_mem[20850] = 0;
disk_mem[20851] = 0;
disk_mem[20852] = 0;
disk_mem[20853] = 0;
disk_mem[20854] = 0;
disk_mem[20855] = 0;
disk_mem[20856] = 0;
disk_mem[20857] = 0;
disk_mem[20858] = 0;
disk_mem[20859] = 0;
disk_mem[20860] = 0;
disk_mem[20861] = 0;
disk_mem[20862] = 0;
disk_mem[20863] = 0;
disk_mem[20864] = 0;
disk_mem[20865] = 0;
disk_mem[20866] = 0;
disk_mem[20867] = 0;
disk_mem[20868] = 0;
disk_mem[20869] = 0;
disk_mem[20870] = 0;
disk_mem[20871] = 0;
disk_mem[20872] = 0;
disk_mem[20873] = 0;
disk_mem[20874] = 0;
disk_mem[20875] = 0;
disk_mem[20876] = 0;
disk_mem[20877] = 0;
disk_mem[20878] = 0;
disk_mem[20879] = 0;
disk_mem[20880] = 0;
disk_mem[20881] = 0;
disk_mem[20882] = 0;
disk_mem[20883] = 0;
disk_mem[20884] = 0;
disk_mem[20885] = 0;
disk_mem[20886] = 0;
disk_mem[20887] = 0;
disk_mem[20888] = 0;
disk_mem[20889] = 0;
disk_mem[20890] = 0;
disk_mem[20891] = 0;
disk_mem[20892] = 0;
disk_mem[20893] = 0;
disk_mem[20894] = 0;
disk_mem[20895] = 0;
disk_mem[20896] = 0;
disk_mem[20897] = 0;
disk_mem[20898] = 0;
disk_mem[20899] = 0;
disk_mem[20900] = 0;
disk_mem[20901] = 0;
disk_mem[20902] = 0;
disk_mem[20903] = 0;
disk_mem[20904] = 0;
disk_mem[20905] = 0;
disk_mem[20906] = 0;
disk_mem[20907] = 0;
disk_mem[20908] = 0;
disk_mem[20909] = 0;
disk_mem[20910] = 0;
disk_mem[20911] = 0;
disk_mem[20912] = 0;
disk_mem[20913] = 0;
disk_mem[20914] = 0;
disk_mem[20915] = 0;
disk_mem[20916] = 0;
disk_mem[20917] = 0;
disk_mem[20918] = 0;
disk_mem[20919] = 0;
disk_mem[20920] = 0;
disk_mem[20921] = 0;
disk_mem[20922] = 0;
disk_mem[20923] = 0;
disk_mem[20924] = 0;
disk_mem[20925] = 0;
disk_mem[20926] = 0;
disk_mem[20927] = 0;
disk_mem[20928] = 0;
disk_mem[20929] = 0;
disk_mem[20930] = 0;
disk_mem[20931] = 0;
disk_mem[20932] = 0;
disk_mem[20933] = 0;
disk_mem[20934] = 0;
disk_mem[20935] = 0;
disk_mem[20936] = 0;
disk_mem[20937] = 0;
disk_mem[20938] = 0;
disk_mem[20939] = 0;
disk_mem[20940] = 0;
disk_mem[20941] = 0;
disk_mem[20942] = 0;
disk_mem[20943] = 0;
disk_mem[20944] = 0;
disk_mem[20945] = 0;
disk_mem[20946] = 0;
disk_mem[20947] = 0;
disk_mem[20948] = 0;
disk_mem[20949] = 0;
disk_mem[20950] = 0;
disk_mem[20951] = 0;
disk_mem[20952] = 0;
disk_mem[20953] = 0;
disk_mem[20954] = 0;
disk_mem[20955] = 0;
disk_mem[20956] = 0;
disk_mem[20957] = 0;
disk_mem[20958] = 0;
disk_mem[20959] = 0;
disk_mem[20960] = 0;
disk_mem[20961] = 0;
disk_mem[20962] = 0;
disk_mem[20963] = 0;
disk_mem[20964] = 0;
disk_mem[20965] = 0;
disk_mem[20966] = 0;
disk_mem[20967] = 0;
disk_mem[20968] = 0;
disk_mem[20969] = 0;
disk_mem[20970] = 0;
disk_mem[20971] = 0;
disk_mem[20972] = 0;
disk_mem[20973] = 0;
disk_mem[20974] = 0;
disk_mem[20975] = 0;
disk_mem[20976] = 0;
disk_mem[20977] = 0;
disk_mem[20978] = 0;
disk_mem[20979] = 0;
disk_mem[20980] = 0;
disk_mem[20981] = 0;
disk_mem[20982] = 0;
disk_mem[20983] = 0;
disk_mem[20984] = 0;
disk_mem[20985] = 0;
disk_mem[20986] = 0;
disk_mem[20987] = 0;
disk_mem[20988] = 0;
disk_mem[20989] = 0;
disk_mem[20990] = 0;
disk_mem[20991] = 0;
disk_mem[20992] = 'h2E;
disk_mem[20993] = 'h20;
disk_mem[20994] = 'h20;
disk_mem[20995] = 'h20;
disk_mem[20996] = 'h20;
disk_mem[20997] = 'h20;
disk_mem[20998] = 'h20;
disk_mem[20999] = 'h20;
disk_mem[21000] = 'h20;
disk_mem[21001] = 'h20;
disk_mem[21002] = 'h20;
disk_mem[21003] = 'h10;
disk_mem[21004] = 0;
disk_mem[21005] = 'h8B;
disk_mem[21006] = 'h90;
disk_mem[21007] = 'h80;
disk_mem[21008] = 'h43;
disk_mem[21009] = 'h55;
disk_mem[21010] = 'h43;
disk_mem[21011] = 'h55;
disk_mem[21012] = 0;
disk_mem[21013] = 0;
disk_mem[21014] = 'h91;
disk_mem[21015] = 'h80;
disk_mem[21016] = 'h43;
disk_mem[21017] = 'h55;
disk_mem[21018] = 'h02;
disk_mem[21019] = 0;
disk_mem[21020] = 0;
disk_mem[21021] = 0;
disk_mem[21022] = 0;
disk_mem[21023] = 0;
disk_mem[21024] = 'h2E;
disk_mem[21025] = 'h2E;
disk_mem[21026] = 'h20;
disk_mem[21027] = 'h20;
disk_mem[21028] = 'h20;
disk_mem[21029] = 'h20;
disk_mem[21030] = 'h20;
disk_mem[21031] = 'h20;
disk_mem[21032] = 'h20;
disk_mem[21033] = 'h20;
disk_mem[21034] = 'h20;
disk_mem[21035] = 'h10;
disk_mem[21036] = 0;
disk_mem[21037] = 'h8B;
disk_mem[21038] = 'h90;
disk_mem[21039] = 'h80;
disk_mem[21040] = 'h43;
disk_mem[21041] = 'h55;
disk_mem[21042] = 'h43;
disk_mem[21043] = 'h55;
disk_mem[21044] = 0;
disk_mem[21045] = 0;
disk_mem[21046] = 'h91;
disk_mem[21047] = 'h80;
disk_mem[21048] = 'h43;
disk_mem[21049] = 'h55;
disk_mem[21050] = 0;
disk_mem[21051] = 0;
disk_mem[21052] = 0;
disk_mem[21053] = 0;
disk_mem[21054] = 0;
disk_mem[21055] = 0;
disk_mem[21056] = 'h42;
disk_mem[21057] = 'h74;
disk_mem[21058] = 0;
disk_mem[21059] = 0;
disk_mem[21060] = 0;
disk_mem[21061] = 'hFF;
disk_mem[21062] = 'hFF;
disk_mem[21063] = 'hFF;
disk_mem[21064] = 'hFF;
disk_mem[21065] = 'hFF;
disk_mem[21066] = 'hFF;
disk_mem[21067] = 'h0F;
disk_mem[21068] = 0;
disk_mem[21069] = 'hCE;
disk_mem[21070] = 'hFF;
disk_mem[21071] = 'hFF;
disk_mem[21072] = 'hFF;
disk_mem[21073] = 'hFF;
disk_mem[21074] = 'hFF;
disk_mem[21075] = 'hFF;
disk_mem[21076] = 'hFF;
disk_mem[21077] = 'hFF;
disk_mem[21078] = 'hFF;
disk_mem[21079] = 'hFF;
disk_mem[21080] = 'hFF;
disk_mem[21081] = 'hFF;
disk_mem[21082] = 0;
disk_mem[21083] = 0;
disk_mem[21084] = 'hFF;
disk_mem[21085] = 'hFF;
disk_mem[21086] = 'hFF;
disk_mem[21087] = 'hFF;
disk_mem[21088] = 'h01;
disk_mem[21089] = 'h57;
disk_mem[21090] = 0;
disk_mem[21091] = 'h50;
disk_mem[21092] = 0;
disk_mem[21093] = 'h53;
disk_mem[21094] = 0;
disk_mem[21095] = 'h65;
disk_mem[21096] = 0;
disk_mem[21097] = 'h74;
disk_mem[21098] = 0;
disk_mem[21099] = 'h0F;
disk_mem[21100] = 0;
disk_mem[21101] = 'hCE;
disk_mem[21102] = 'h74;
disk_mem[21103] = 0;
disk_mem[21104] = 'h69;
disk_mem[21105] = 0;
disk_mem[21106] = 'h6E;
disk_mem[21107] = 0;
disk_mem[21108] = 'h67;
disk_mem[21109] = 0;
disk_mem[21110] = 'h73;
disk_mem[21111] = 0;
disk_mem[21112] = 'h2E;
disk_mem[21113] = 0;
disk_mem[21114] = 0;
disk_mem[21115] = 0;
disk_mem[21116] = 'h64;
disk_mem[21117] = 0;
disk_mem[21118] = 'h61;
disk_mem[21119] = 0;
disk_mem[21120] = 'h57;
disk_mem[21121] = 'h50;
disk_mem[21122] = 'h53;
disk_mem[21123] = 'h45;
disk_mem[21124] = 'h54;
disk_mem[21125] = 'h54;
disk_mem[21126] = 'h7E;
disk_mem[21127] = 'h31;
disk_mem[21128] = 'h44;
disk_mem[21129] = 'h41;
disk_mem[21130] = 'h54;
disk_mem[21131] = 'h20;
disk_mem[21132] = 0;
disk_mem[21133] = 'h93;
disk_mem[21134] = 'h90;
disk_mem[21135] = 'h80;
disk_mem[21136] = 'h43;
disk_mem[21137] = 'h55;
disk_mem[21138] = 'h43;
disk_mem[21139] = 'h55;
disk_mem[21140] = 0;
disk_mem[21141] = 0;
disk_mem[21142] = 'h91;
disk_mem[21143] = 'h80;
disk_mem[21144] = 'h43;
disk_mem[21145] = 'h55;
disk_mem[21146] = 'h03;
disk_mem[21147] = 0;
disk_mem[21148] = 'h0C;
disk_mem[21149] = 0;
disk_mem[21150] = 0;
disk_mem[21151] = 0;
disk_mem[21152] = 'h42;
disk_mem[21153] = 'h47;
disk_mem[21154] = 0;
disk_mem[21155] = 'h75;
disk_mem[21156] = 0;
disk_mem[21157] = 'h69;
disk_mem[21158] = 0;
disk_mem[21159] = 'h64;
disk_mem[21160] = 0;
disk_mem[21161] = 0;
disk_mem[21162] = 0;
disk_mem[21163] = 'h0F;
disk_mem[21164] = 0;
disk_mem[21165] = 'hFF;
disk_mem[21166] = 'hFF;
disk_mem[21167] = 'hFF;
disk_mem[21168] = 'hFF;
disk_mem[21169] = 'hFF;
disk_mem[21170] = 'hFF;
disk_mem[21171] = 'hFF;
disk_mem[21172] = 'hFF;
disk_mem[21173] = 'hFF;
disk_mem[21174] = 'hFF;
disk_mem[21175] = 'hFF;
disk_mem[21176] = 'hFF;
disk_mem[21177] = 'hFF;
disk_mem[21178] = 0;
disk_mem[21179] = 0;
disk_mem[21180] = 'hFF;
disk_mem[21181] = 'hFF;
disk_mem[21182] = 'hFF;
disk_mem[21183] = 'hFF;
disk_mem[21184] = 'h01;
disk_mem[21185] = 'h49;
disk_mem[21186] = 0;
disk_mem[21187] = 'h6E;
disk_mem[21188] = 0;
disk_mem[21189] = 'h64;
disk_mem[21190] = 0;
disk_mem[21191] = 'h65;
disk_mem[21192] = 0;
disk_mem[21193] = 'h78;
disk_mem[21194] = 0;
disk_mem[21195] = 'h0F;
disk_mem[21196] = 0;
disk_mem[21197] = 'hFF;
disk_mem[21198] = 'h65;
disk_mem[21199] = 0;
disk_mem[21200] = 'h72;
disk_mem[21201] = 0;
disk_mem[21202] = 'h56;
disk_mem[21203] = 0;
disk_mem[21204] = 'h6F;
disk_mem[21205] = 0;
disk_mem[21206] = 'h6C;
disk_mem[21207] = 0;
disk_mem[21208] = 'h75;
disk_mem[21209] = 0;
disk_mem[21210] = 0;
disk_mem[21211] = 0;
disk_mem[21212] = 'h6D;
disk_mem[21213] = 0;
disk_mem[21214] = 'h65;
disk_mem[21215] = 0;
disk_mem[21216] = 'h49;
disk_mem[21217] = 'h4E;
disk_mem[21218] = 'h44;
disk_mem[21219] = 'h45;
disk_mem[21220] = 'h58;
disk_mem[21221] = 'h45;
disk_mem[21222] = 'h7E;
disk_mem[21223] = 'h31;
disk_mem[21224] = 'h20;
disk_mem[21225] = 'h20;
disk_mem[21226] = 'h20;
disk_mem[21227] = 'h20;
disk_mem[21228] = 0;
disk_mem[21229] = 'h22;
disk_mem[21230] = 'h93;
disk_mem[21231] = 'h80;
disk_mem[21232] = 'h43;
disk_mem[21233] = 'h55;
disk_mem[21234] = 'h43;
disk_mem[21235] = 'h55;
disk_mem[21236] = 0;
disk_mem[21237] = 0;
disk_mem[21238] = 'h94;
disk_mem[21239] = 'h80;
disk_mem[21240] = 'h43;
disk_mem[21241] = 'h55;
disk_mem[21242] = 'h04;
disk_mem[21243] = 0;
disk_mem[21244] = 'h4C;
disk_mem[21245] = 0;
disk_mem[21246] = 0;
disk_mem[21247] = 0;
disk_mem[21248] = 0;
disk_mem[21249] = 0;
disk_mem[21250] = 0;
disk_mem[21251] = 0;
disk_mem[21252] = 0;
disk_mem[21253] = 0;
disk_mem[21254] = 0;
disk_mem[21255] = 0;
disk_mem[21256] = 0;
disk_mem[21257] = 0;
disk_mem[21258] = 0;
disk_mem[21259] = 0;
disk_mem[21260] = 0;
disk_mem[21261] = 0;
disk_mem[21262] = 0;
disk_mem[21263] = 0;
disk_mem[21264] = 0;
disk_mem[21265] = 0;
disk_mem[21266] = 0;
disk_mem[21267] = 0;
disk_mem[21268] = 0;
disk_mem[21269] = 0;
disk_mem[21270] = 0;
disk_mem[21271] = 0;
disk_mem[21272] = 0;
disk_mem[21273] = 0;
disk_mem[21274] = 0;
disk_mem[21275] = 0;
disk_mem[21276] = 0;
disk_mem[21277] = 0;
disk_mem[21278] = 0;
disk_mem[21279] = 0;
disk_mem[21280] = 0;
disk_mem[21281] = 0;
disk_mem[21282] = 0;
disk_mem[21283] = 0;
disk_mem[21284] = 0;
disk_mem[21285] = 0;
disk_mem[21286] = 0;
disk_mem[21287] = 0;
disk_mem[21288] = 0;
disk_mem[21289] = 0;
disk_mem[21290] = 0;
disk_mem[21291] = 0;
disk_mem[21292] = 0;
disk_mem[21293] = 0;
disk_mem[21294] = 0;
disk_mem[21295] = 0;
disk_mem[21296] = 0;
disk_mem[21297] = 0;
disk_mem[21298] = 0;
disk_mem[21299] = 0;
disk_mem[21300] = 0;
disk_mem[21301] = 0;
disk_mem[21302] = 0;
disk_mem[21303] = 0;
disk_mem[21304] = 0;
disk_mem[21305] = 0;
disk_mem[21306] = 0;
disk_mem[21307] = 0;
disk_mem[21308] = 0;
disk_mem[21309] = 0;
disk_mem[21310] = 0;
disk_mem[21311] = 0;
disk_mem[21312] = 0;
disk_mem[21313] = 0;
disk_mem[21314] = 0;
disk_mem[21315] = 0;
disk_mem[21316] = 0;
disk_mem[21317] = 0;
disk_mem[21318] = 0;
disk_mem[21319] = 0;
disk_mem[21320] = 0;
disk_mem[21321] = 0;
disk_mem[21322] = 0;
disk_mem[21323] = 0;
disk_mem[21324] = 0;
disk_mem[21325] = 0;
disk_mem[21326] = 0;
disk_mem[21327] = 0;
disk_mem[21328] = 0;
disk_mem[21329] = 0;
disk_mem[21330] = 0;
disk_mem[21331] = 0;
disk_mem[21332] = 0;
disk_mem[21333] = 0;
disk_mem[21334] = 0;
disk_mem[21335] = 0;
disk_mem[21336] = 0;
disk_mem[21337] = 0;
disk_mem[21338] = 0;
disk_mem[21339] = 0;
disk_mem[21340] = 0;
disk_mem[21341] = 0;
disk_mem[21342] = 0;
disk_mem[21343] = 0;
disk_mem[21344] = 0;
disk_mem[21345] = 0;
disk_mem[21346] = 0;
disk_mem[21347] = 0;
disk_mem[21348] = 0;
disk_mem[21349] = 0;
disk_mem[21350] = 0;
disk_mem[21351] = 0;
disk_mem[21352] = 0;
disk_mem[21353] = 0;
disk_mem[21354] = 0;
disk_mem[21355] = 0;
disk_mem[21356] = 0;
disk_mem[21357] = 0;
disk_mem[21358] = 0;
disk_mem[21359] = 0;
disk_mem[21360] = 0;
disk_mem[21361] = 0;
disk_mem[21362] = 0;
disk_mem[21363] = 0;
disk_mem[21364] = 0;
disk_mem[21365] = 0;
disk_mem[21366] = 0;
disk_mem[21367] = 0;
disk_mem[21368] = 0;
disk_mem[21369] = 0;
disk_mem[21370] = 0;
disk_mem[21371] = 0;
disk_mem[21372] = 0;
disk_mem[21373] = 0;
disk_mem[21374] = 0;
disk_mem[21375] = 0;
disk_mem[21376] = 0;
disk_mem[21377] = 0;
disk_mem[21378] = 0;
disk_mem[21379] = 0;
disk_mem[21380] = 0;
disk_mem[21381] = 0;
disk_mem[21382] = 0;
disk_mem[21383] = 0;
disk_mem[21384] = 0;
disk_mem[21385] = 0;
disk_mem[21386] = 0;
disk_mem[21387] = 0;
disk_mem[21388] = 0;
disk_mem[21389] = 0;
disk_mem[21390] = 0;
disk_mem[21391] = 0;
disk_mem[21392] = 0;
disk_mem[21393] = 0;
disk_mem[21394] = 0;
disk_mem[21395] = 0;
disk_mem[21396] = 0;
disk_mem[21397] = 0;
disk_mem[21398] = 0;
disk_mem[21399] = 0;
disk_mem[21400] = 0;
disk_mem[21401] = 0;
disk_mem[21402] = 0;
disk_mem[21403] = 0;
disk_mem[21404] = 0;
disk_mem[21405] = 0;
disk_mem[21406] = 0;
disk_mem[21407] = 0;
disk_mem[21408] = 0;
disk_mem[21409] = 0;
disk_mem[21410] = 0;
disk_mem[21411] = 0;
disk_mem[21412] = 0;
disk_mem[21413] = 0;
disk_mem[21414] = 0;
disk_mem[21415] = 0;
disk_mem[21416] = 0;
disk_mem[21417] = 0;
disk_mem[21418] = 0;
disk_mem[21419] = 0;
disk_mem[21420] = 0;
disk_mem[21421] = 0;
disk_mem[21422] = 0;
disk_mem[21423] = 0;
disk_mem[21424] = 0;
disk_mem[21425] = 0;
disk_mem[21426] = 0;
disk_mem[21427] = 0;
disk_mem[21428] = 0;
disk_mem[21429] = 0;
disk_mem[21430] = 0;
disk_mem[21431] = 0;
disk_mem[21432] = 0;
disk_mem[21433] = 0;
disk_mem[21434] = 0;
disk_mem[21435] = 0;
disk_mem[21436] = 0;
disk_mem[21437] = 0;
disk_mem[21438] = 0;
disk_mem[21439] = 0;
disk_mem[21440] = 0;
disk_mem[21441] = 0;
disk_mem[21442] = 0;
disk_mem[21443] = 0;
disk_mem[21444] = 0;
disk_mem[21445] = 0;
disk_mem[21446] = 0;
disk_mem[21447] = 0;
disk_mem[21448] = 0;
disk_mem[21449] = 0;
disk_mem[21450] = 0;
disk_mem[21451] = 0;
disk_mem[21452] = 0;
disk_mem[21453] = 0;
disk_mem[21454] = 0;
disk_mem[21455] = 0;
disk_mem[21456] = 0;
disk_mem[21457] = 0;
disk_mem[21458] = 0;
disk_mem[21459] = 0;
disk_mem[21460] = 0;
disk_mem[21461] = 0;
disk_mem[21462] = 0;
disk_mem[21463] = 0;
disk_mem[21464] = 0;
disk_mem[21465] = 0;
disk_mem[21466] = 0;
disk_mem[21467] = 0;
disk_mem[21468] = 0;
disk_mem[21469] = 0;
disk_mem[21470] = 0;
disk_mem[21471] = 0;
disk_mem[21472] = 0;
disk_mem[21473] = 0;
disk_mem[21474] = 0;
disk_mem[21475] = 0;
disk_mem[21476] = 0;
disk_mem[21477] = 0;
disk_mem[21478] = 0;
disk_mem[21479] = 0;
disk_mem[21480] = 0;
disk_mem[21481] = 0;
disk_mem[21482] = 0;
disk_mem[21483] = 0;
disk_mem[21484] = 0;
disk_mem[21485] = 0;
disk_mem[21486] = 0;
disk_mem[21487] = 0;
disk_mem[21488] = 0;
disk_mem[21489] = 0;
disk_mem[21490] = 0;
disk_mem[21491] = 0;
disk_mem[21492] = 0;
disk_mem[21493] = 0;
disk_mem[21494] = 0;
disk_mem[21495] = 0;
disk_mem[21496] = 0;
disk_mem[21497] = 0;
disk_mem[21498] = 0;
disk_mem[21499] = 0;
disk_mem[21500] = 0;
disk_mem[21501] = 0;
disk_mem[21502] = 0;
disk_mem[21503] = 0;
disk_mem[21504] = 'h0C;
disk_mem[21505] = 0;
disk_mem[21506] = 0;
disk_mem[21507] = 0;
disk_mem[21508] = 'hED;
disk_mem[21509] = 'hEF;
disk_mem[21510] = 'hF3;
disk_mem[21511] = 'hF7;
disk_mem[21512] = 0;
disk_mem[21513] = 'hEB;
disk_mem[21514] = 'h4F;
disk_mem[21515] = 'hE2;
disk_mem[21516] = 0;
disk_mem[21517] = 0;
disk_mem[21518] = 0;
disk_mem[21519] = 0;
disk_mem[21520] = 0;
disk_mem[21521] = 0;
disk_mem[21522] = 0;
disk_mem[21523] = 0;
disk_mem[21524] = 0;
disk_mem[21525] = 0;
disk_mem[21526] = 0;
disk_mem[21527] = 0;
disk_mem[21528] = 0;
disk_mem[21529] = 0;
disk_mem[21530] = 0;
disk_mem[21531] = 0;
disk_mem[21532] = 0;
disk_mem[21533] = 0;
disk_mem[21534] = 0;
disk_mem[21535] = 0;
disk_mem[21536] = 0;
disk_mem[21537] = 0;
disk_mem[21538] = 0;
disk_mem[21539] = 0;
disk_mem[21540] = 0;
disk_mem[21541] = 0;
disk_mem[21542] = 0;
disk_mem[21543] = 0;
disk_mem[21544] = 0;
disk_mem[21545] = 0;
disk_mem[21546] = 0;
disk_mem[21547] = 0;
disk_mem[21548] = 0;
disk_mem[21549] = 0;
disk_mem[21550] = 0;
disk_mem[21551] = 0;
disk_mem[21552] = 0;
disk_mem[21553] = 0;
disk_mem[21554] = 0;
disk_mem[21555] = 0;
disk_mem[21556] = 0;
disk_mem[21557] = 0;
disk_mem[21558] = 0;
disk_mem[21559] = 0;
disk_mem[21560] = 0;
disk_mem[21561] = 0;
disk_mem[21562] = 0;
disk_mem[21563] = 0;
disk_mem[21564] = 0;
disk_mem[21565] = 0;
disk_mem[21566] = 0;
disk_mem[21567] = 0;
disk_mem[21568] = 0;
disk_mem[21569] = 0;
disk_mem[21570] = 0;
disk_mem[21571] = 0;
disk_mem[21572] = 0;
disk_mem[21573] = 0;
disk_mem[21574] = 0;
disk_mem[21575] = 0;
disk_mem[21576] = 0;
disk_mem[21577] = 0;
disk_mem[21578] = 0;
disk_mem[21579] = 0;
disk_mem[21580] = 0;
disk_mem[21581] = 0;
disk_mem[21582] = 0;
disk_mem[21583] = 0;
disk_mem[21584] = 0;
disk_mem[21585] = 0;
disk_mem[21586] = 0;
disk_mem[21587] = 0;
disk_mem[21588] = 0;
disk_mem[21589] = 0;
disk_mem[21590] = 0;
disk_mem[21591] = 0;
disk_mem[21592] = 0;
disk_mem[21593] = 0;
disk_mem[21594] = 0;
disk_mem[21595] = 0;
disk_mem[21596] = 0;
disk_mem[21597] = 0;
disk_mem[21598] = 0;
disk_mem[21599] = 0;
disk_mem[21600] = 0;
disk_mem[21601] = 0;
disk_mem[21602] = 0;
disk_mem[21603] = 0;
disk_mem[21604] = 0;
disk_mem[21605] = 0;
disk_mem[21606] = 0;
disk_mem[21607] = 0;
disk_mem[21608] = 0;
disk_mem[21609] = 0;
disk_mem[21610] = 0;
disk_mem[21611] = 0;
disk_mem[21612] = 0;
disk_mem[21613] = 0;
disk_mem[21614] = 0;
disk_mem[21615] = 0;
disk_mem[21616] = 0;
disk_mem[21617] = 0;
disk_mem[21618] = 0;
disk_mem[21619] = 0;
disk_mem[21620] = 0;
disk_mem[21621] = 0;
disk_mem[21622] = 0;
disk_mem[21623] = 0;
disk_mem[21624] = 0;
disk_mem[21625] = 0;
disk_mem[21626] = 0;
disk_mem[21627] = 0;
disk_mem[21628] = 0;
disk_mem[21629] = 0;
disk_mem[21630] = 0;
disk_mem[21631] = 0;
disk_mem[21632] = 0;
disk_mem[21633] = 0;
disk_mem[21634] = 0;
disk_mem[21635] = 0;
disk_mem[21636] = 0;
disk_mem[21637] = 0;
disk_mem[21638] = 0;
disk_mem[21639] = 0;
disk_mem[21640] = 0;
disk_mem[21641] = 0;
disk_mem[21642] = 0;
disk_mem[21643] = 0;
disk_mem[21644] = 0;
disk_mem[21645] = 0;
disk_mem[21646] = 0;
disk_mem[21647] = 0;
disk_mem[21648] = 0;
disk_mem[21649] = 0;
disk_mem[21650] = 0;
disk_mem[21651] = 0;
disk_mem[21652] = 0;
disk_mem[21653] = 0;
disk_mem[21654] = 0;
disk_mem[21655] = 0;
disk_mem[21656] = 0;
disk_mem[21657] = 0;
disk_mem[21658] = 0;
disk_mem[21659] = 0;
disk_mem[21660] = 0;
disk_mem[21661] = 0;
disk_mem[21662] = 0;
disk_mem[21663] = 0;
disk_mem[21664] = 0;
disk_mem[21665] = 0;
disk_mem[21666] = 0;
disk_mem[21667] = 0;
disk_mem[21668] = 0;
disk_mem[21669] = 0;
disk_mem[21670] = 0;
disk_mem[21671] = 0;
disk_mem[21672] = 0;
disk_mem[21673] = 0;
disk_mem[21674] = 0;
disk_mem[21675] = 0;
disk_mem[21676] = 0;
disk_mem[21677] = 0;
disk_mem[21678] = 0;
disk_mem[21679] = 0;
disk_mem[21680] = 0;
disk_mem[21681] = 0;
disk_mem[21682] = 0;
disk_mem[21683] = 0;
disk_mem[21684] = 0;
disk_mem[21685] = 0;
disk_mem[21686] = 0;
disk_mem[21687] = 0;
disk_mem[21688] = 0;
disk_mem[21689] = 0;
disk_mem[21690] = 0;
disk_mem[21691] = 0;
disk_mem[21692] = 0;
disk_mem[21693] = 0;
disk_mem[21694] = 0;
disk_mem[21695] = 0;
disk_mem[21696] = 0;
disk_mem[21697] = 0;
disk_mem[21698] = 0;
disk_mem[21699] = 0;
disk_mem[21700] = 0;
disk_mem[21701] = 0;
disk_mem[21702] = 0;
disk_mem[21703] = 0;
disk_mem[21704] = 0;
disk_mem[21705] = 0;
disk_mem[21706] = 0;
disk_mem[21707] = 0;
disk_mem[21708] = 0;
disk_mem[21709] = 0;
disk_mem[21710] = 0;
disk_mem[21711] = 0;
disk_mem[21712] = 0;
disk_mem[21713] = 0;
disk_mem[21714] = 0;
disk_mem[21715] = 0;
disk_mem[21716] = 0;
disk_mem[21717] = 0;
disk_mem[21718] = 0;
disk_mem[21719] = 0;
disk_mem[21720] = 0;
disk_mem[21721] = 0;
disk_mem[21722] = 0;
disk_mem[21723] = 0;
disk_mem[21724] = 0;
disk_mem[21725] = 0;
disk_mem[21726] = 0;
disk_mem[21727] = 0;
disk_mem[21728] = 0;
disk_mem[21729] = 0;
disk_mem[21730] = 0;
disk_mem[21731] = 0;
disk_mem[21732] = 0;
disk_mem[21733] = 0;
disk_mem[21734] = 0;
disk_mem[21735] = 0;
disk_mem[21736] = 0;
disk_mem[21737] = 0;
disk_mem[21738] = 0;
disk_mem[21739] = 0;
disk_mem[21740] = 0;
disk_mem[21741] = 0;
disk_mem[21742] = 0;
disk_mem[21743] = 0;
disk_mem[21744] = 0;
disk_mem[21745] = 0;
disk_mem[21746] = 0;
disk_mem[21747] = 0;
disk_mem[21748] = 0;
disk_mem[21749] = 0;
disk_mem[21750] = 0;
disk_mem[21751] = 0;
disk_mem[21752] = 0;
disk_mem[21753] = 0;
disk_mem[21754] = 0;
disk_mem[21755] = 0;
disk_mem[21756] = 0;
disk_mem[21757] = 0;
disk_mem[21758] = 0;
disk_mem[21759] = 0;
disk_mem[21760] = 0;
disk_mem[21761] = 0;
disk_mem[21762] = 0;
disk_mem[21763] = 0;
disk_mem[21764] = 0;
disk_mem[21765] = 0;
disk_mem[21766] = 0;
disk_mem[21767] = 0;
disk_mem[21768] = 0;
disk_mem[21769] = 0;
disk_mem[21770] = 0;
disk_mem[21771] = 0;
disk_mem[21772] = 0;
disk_mem[21773] = 0;
disk_mem[21774] = 0;
disk_mem[21775] = 0;
disk_mem[21776] = 0;
disk_mem[21777] = 0;
disk_mem[21778] = 0;
disk_mem[21779] = 0;
disk_mem[21780] = 0;
disk_mem[21781] = 0;
disk_mem[21782] = 0;
disk_mem[21783] = 0;
disk_mem[21784] = 0;
disk_mem[21785] = 0;
disk_mem[21786] = 0;
disk_mem[21787] = 0;
disk_mem[21788] = 0;
disk_mem[21789] = 0;
disk_mem[21790] = 0;
disk_mem[21791] = 0;
disk_mem[21792] = 0;
disk_mem[21793] = 0;
disk_mem[21794] = 0;
disk_mem[21795] = 0;
disk_mem[21796] = 0;
disk_mem[21797] = 0;
disk_mem[21798] = 0;
disk_mem[21799] = 0;
disk_mem[21800] = 0;
disk_mem[21801] = 0;
disk_mem[21802] = 0;
disk_mem[21803] = 0;
disk_mem[21804] = 0;
disk_mem[21805] = 0;
disk_mem[21806] = 0;
disk_mem[21807] = 0;
disk_mem[21808] = 0;
disk_mem[21809] = 0;
disk_mem[21810] = 0;
disk_mem[21811] = 0;
disk_mem[21812] = 0;
disk_mem[21813] = 0;
disk_mem[21814] = 0;
disk_mem[21815] = 0;
disk_mem[21816] = 0;
disk_mem[21817] = 0;
disk_mem[21818] = 0;
disk_mem[21819] = 0;
disk_mem[21820] = 0;
disk_mem[21821] = 0;
disk_mem[21822] = 0;
disk_mem[21823] = 0;
disk_mem[21824] = 0;
disk_mem[21825] = 0;
disk_mem[21826] = 0;
disk_mem[21827] = 0;
disk_mem[21828] = 0;
disk_mem[21829] = 0;
disk_mem[21830] = 0;
disk_mem[21831] = 0;
disk_mem[21832] = 0;
disk_mem[21833] = 0;
disk_mem[21834] = 0;
disk_mem[21835] = 0;
disk_mem[21836] = 0;
disk_mem[21837] = 0;
disk_mem[21838] = 0;
disk_mem[21839] = 0;
disk_mem[21840] = 0;
disk_mem[21841] = 0;
disk_mem[21842] = 0;
disk_mem[21843] = 0;
disk_mem[21844] = 0;
disk_mem[21845] = 0;
disk_mem[21846] = 0;
disk_mem[21847] = 0;
disk_mem[21848] = 0;
disk_mem[21849] = 0;
disk_mem[21850] = 0;
disk_mem[21851] = 0;
disk_mem[21852] = 0;
disk_mem[21853] = 0;
disk_mem[21854] = 0;
disk_mem[21855] = 0;
disk_mem[21856] = 0;
disk_mem[21857] = 0;
disk_mem[21858] = 0;
disk_mem[21859] = 0;
disk_mem[21860] = 0;
disk_mem[21861] = 0;
disk_mem[21862] = 0;
disk_mem[21863] = 0;
disk_mem[21864] = 0;
disk_mem[21865] = 0;
disk_mem[21866] = 0;
disk_mem[21867] = 0;
disk_mem[21868] = 0;
disk_mem[21869] = 0;
disk_mem[21870] = 0;
disk_mem[21871] = 0;
disk_mem[21872] = 0;
disk_mem[21873] = 0;
disk_mem[21874] = 0;
disk_mem[21875] = 0;
disk_mem[21876] = 0;
disk_mem[21877] = 0;
disk_mem[21878] = 0;
disk_mem[21879] = 0;
disk_mem[21880] = 0;
disk_mem[21881] = 0;
disk_mem[21882] = 0;
disk_mem[21883] = 0;
disk_mem[21884] = 0;
disk_mem[21885] = 0;
disk_mem[21886] = 0;
disk_mem[21887] = 0;
disk_mem[21888] = 0;
disk_mem[21889] = 0;
disk_mem[21890] = 0;
disk_mem[21891] = 0;
disk_mem[21892] = 0;
disk_mem[21893] = 0;
disk_mem[21894] = 0;
disk_mem[21895] = 0;
disk_mem[21896] = 0;
disk_mem[21897] = 0;
disk_mem[21898] = 0;
disk_mem[21899] = 0;
disk_mem[21900] = 0;
disk_mem[21901] = 0;
disk_mem[21902] = 0;
disk_mem[21903] = 0;
disk_mem[21904] = 0;
disk_mem[21905] = 0;
disk_mem[21906] = 0;
disk_mem[21907] = 0;
disk_mem[21908] = 0;
disk_mem[21909] = 0;
disk_mem[21910] = 0;
disk_mem[21911] = 0;
disk_mem[21912] = 0;
disk_mem[21913] = 0;
disk_mem[21914] = 0;
disk_mem[21915] = 0;
disk_mem[21916] = 0;
disk_mem[21917] = 0;
disk_mem[21918] = 0;
disk_mem[21919] = 0;
disk_mem[21920] = 0;
disk_mem[21921] = 0;
disk_mem[21922] = 0;
disk_mem[21923] = 0;
disk_mem[21924] = 0;
disk_mem[21925] = 0;
disk_mem[21926] = 0;
disk_mem[21927] = 0;
disk_mem[21928] = 0;
disk_mem[21929] = 0;
disk_mem[21930] = 0;
disk_mem[21931] = 0;
disk_mem[21932] = 0;
disk_mem[21933] = 0;
disk_mem[21934] = 0;
disk_mem[21935] = 0;
disk_mem[21936] = 0;
disk_mem[21937] = 0;
disk_mem[21938] = 0;
disk_mem[21939] = 0;
disk_mem[21940] = 0;
disk_mem[21941] = 0;
disk_mem[21942] = 0;
disk_mem[21943] = 0;
disk_mem[21944] = 0;
disk_mem[21945] = 0;
disk_mem[21946] = 0;
disk_mem[21947] = 0;
disk_mem[21948] = 0;
disk_mem[21949] = 0;
disk_mem[21950] = 0;
disk_mem[21951] = 0;
disk_mem[21952] = 0;
disk_mem[21953] = 0;
disk_mem[21954] = 0;
disk_mem[21955] = 0;
disk_mem[21956] = 0;
disk_mem[21957] = 0;
disk_mem[21958] = 0;
disk_mem[21959] = 0;
disk_mem[21960] = 0;
disk_mem[21961] = 0;
disk_mem[21962] = 0;
disk_mem[21963] = 0;
disk_mem[21964] = 0;
disk_mem[21965] = 0;
disk_mem[21966] = 0;
disk_mem[21967] = 0;
disk_mem[21968] = 0;
disk_mem[21969] = 0;
disk_mem[21970] = 0;
disk_mem[21971] = 0;
disk_mem[21972] = 0;
disk_mem[21973] = 0;
disk_mem[21974] = 0;
disk_mem[21975] = 0;
disk_mem[21976] = 0;
disk_mem[21977] = 0;
disk_mem[21978] = 0;
disk_mem[21979] = 0;
disk_mem[21980] = 0;
disk_mem[21981] = 0;
disk_mem[21982] = 0;
disk_mem[21983] = 0;
disk_mem[21984] = 0;
disk_mem[21985] = 0;
disk_mem[21986] = 0;
disk_mem[21987] = 0;
disk_mem[21988] = 0;
disk_mem[21989] = 0;
disk_mem[21990] = 0;
disk_mem[21991] = 0;
disk_mem[21992] = 0;
disk_mem[21993] = 0;
disk_mem[21994] = 0;
disk_mem[21995] = 0;
disk_mem[21996] = 0;
disk_mem[21997] = 0;
disk_mem[21998] = 0;
disk_mem[21999] = 0;
disk_mem[22000] = 0;
disk_mem[22001] = 0;
disk_mem[22002] = 0;
disk_mem[22003] = 0;
disk_mem[22004] = 0;
disk_mem[22005] = 0;
disk_mem[22006] = 0;
disk_mem[22007] = 0;
disk_mem[22008] = 0;
disk_mem[22009] = 0;
disk_mem[22010] = 0;
disk_mem[22011] = 0;
disk_mem[22012] = 0;
disk_mem[22013] = 0;
disk_mem[22014] = 0;
disk_mem[22015] = 0;
disk_mem[22016] = 'h7B;
disk_mem[22017] = 0;
disk_mem[22018] = 'h46;
disk_mem[22019] = 0;
disk_mem[22020] = 'h30;
disk_mem[22021] = 0;
disk_mem[22022] = 'h33;
disk_mem[22023] = 0;
disk_mem[22024] = 'h32;
disk_mem[22025] = 0;
disk_mem[22026] = 'h43;
disk_mem[22027] = 0;
disk_mem[22028] = 'h41;
disk_mem[22029] = 0;
disk_mem[22030] = 'h33;
disk_mem[22031] = 0;
disk_mem[22032] = 'h35;
disk_mem[22033] = 0;
disk_mem[22034] = 'h2D;
disk_mem[22035] = 0;
disk_mem[22036] = 'h45;
disk_mem[22037] = 0;
disk_mem[22038] = 'h45;
disk_mem[22039] = 0;
disk_mem[22040] = 'h46;
disk_mem[22041] = 0;
disk_mem[22042] = 'h31;
disk_mem[22043] = 0;
disk_mem[22044] = 'h2D;
disk_mem[22045] = 0;
disk_mem[22046] = 'h34;
disk_mem[22047] = 0;
disk_mem[22048] = 'h35;
disk_mem[22049] = 0;
disk_mem[22050] = 'h44;
disk_mem[22051] = 0;
disk_mem[22052] = 'h30;
disk_mem[22053] = 0;
disk_mem[22054] = 'h2D;
disk_mem[22055] = 0;
disk_mem[22056] = 'h42;
disk_mem[22057] = 0;
disk_mem[22058] = 'h34;
disk_mem[22059] = 0;
disk_mem[22060] = 'h32;
disk_mem[22061] = 0;
disk_mem[22062] = 'h33;
disk_mem[22063] = 0;
disk_mem[22064] = 'h2D;
disk_mem[22065] = 0;
disk_mem[22066] = 'h41;
disk_mem[22067] = 0;
disk_mem[22068] = 'h43;
disk_mem[22069] = 0;
disk_mem[22070] = 'h43;
disk_mem[22071] = 0;
disk_mem[22072] = 'h34;
disk_mem[22073] = 0;
disk_mem[22074] = 'h43;
disk_mem[22075] = 0;
disk_mem[22076] = 'h36;
disk_mem[22077] = 0;
disk_mem[22078] = 'h30;
disk_mem[22079] = 0;
disk_mem[22080] = 'h39;
disk_mem[22081] = 0;
disk_mem[22082] = 'h38;
disk_mem[22083] = 0;
disk_mem[22084] = 'h36;
disk_mem[22085] = 0;
disk_mem[22086] = 'h45;
disk_mem[22087] = 0;
disk_mem[22088] = 'h45;
disk_mem[22089] = 0;
disk_mem[22090] = 'h7D;
disk_mem[22091] = 0;
disk_mem[22092] = 0;
disk_mem[22093] = 0;
disk_mem[22094] = 0;
disk_mem[22095] = 0;
disk_mem[22096] = 0;
disk_mem[22097] = 0;
disk_mem[22098] = 0;
disk_mem[22099] = 0;
disk_mem[22100] = 0;
disk_mem[22101] = 0;
disk_mem[22102] = 0;
disk_mem[22103] = 0;
disk_mem[22104] = 0;
disk_mem[22105] = 0;
disk_mem[22106] = 0;
disk_mem[22107] = 0;
disk_mem[22108] = 0;
disk_mem[22109] = 0;
disk_mem[22110] = 0;
disk_mem[22111] = 0;
disk_mem[22112] = 0;
disk_mem[22113] = 0;
disk_mem[22114] = 0;
disk_mem[22115] = 0;
disk_mem[22116] = 0;
disk_mem[22117] = 0;
disk_mem[22118] = 0;
disk_mem[22119] = 0;
disk_mem[22120] = 0;
disk_mem[22121] = 0;
disk_mem[22122] = 0;
disk_mem[22123] = 0;
disk_mem[22124] = 0;
disk_mem[22125] = 0;
disk_mem[22126] = 0;
disk_mem[22127] = 0;
disk_mem[22128] = 0;
disk_mem[22129] = 0;
disk_mem[22130] = 0;
disk_mem[22131] = 0;
disk_mem[22132] = 0;
disk_mem[22133] = 0;
disk_mem[22134] = 0;
disk_mem[22135] = 0;
disk_mem[22136] = 0;
disk_mem[22137] = 0;
disk_mem[22138] = 0;
disk_mem[22139] = 0;
disk_mem[22140] = 0;
disk_mem[22141] = 0;
disk_mem[22142] = 0;
disk_mem[22143] = 0;
disk_mem[22144] = 0;
disk_mem[22145] = 0;
disk_mem[22146] = 0;
disk_mem[22147] = 0;
disk_mem[22148] = 0;
disk_mem[22149] = 0;
disk_mem[22150] = 0;
disk_mem[22151] = 0;
disk_mem[22152] = 0;
disk_mem[22153] = 0;
disk_mem[22154] = 0;
disk_mem[22155] = 0;
disk_mem[22156] = 0;
disk_mem[22157] = 0;
disk_mem[22158] = 0;
disk_mem[22159] = 0;
disk_mem[22160] = 0;
disk_mem[22161] = 0;
disk_mem[22162] = 0;
disk_mem[22163] = 0;
disk_mem[22164] = 0;
disk_mem[22165] = 0;
disk_mem[22166] = 0;
disk_mem[22167] = 0;
disk_mem[22168] = 0;
disk_mem[22169] = 0;
disk_mem[22170] = 0;
disk_mem[22171] = 0;
disk_mem[22172] = 0;
disk_mem[22173] = 0;
disk_mem[22174] = 0;
disk_mem[22175] = 0;
disk_mem[22176] = 0;
disk_mem[22177] = 0;
disk_mem[22178] = 0;
disk_mem[22179] = 0;
disk_mem[22180] = 0;
disk_mem[22181] = 0;
disk_mem[22182] = 0;
disk_mem[22183] = 0;
disk_mem[22184] = 0;
disk_mem[22185] = 0;
disk_mem[22186] = 0;
disk_mem[22187] = 0;
disk_mem[22188] = 0;
disk_mem[22189] = 0;
disk_mem[22190] = 0;
disk_mem[22191] = 0;
disk_mem[22192] = 0;
disk_mem[22193] = 0;
disk_mem[22194] = 0;
disk_mem[22195] = 0;
disk_mem[22196] = 0;
disk_mem[22197] = 0;
disk_mem[22198] = 0;
disk_mem[22199] = 0;
disk_mem[22200] = 0;
disk_mem[22201] = 0;
disk_mem[22202] = 0;
disk_mem[22203] = 0;
disk_mem[22204] = 0;
disk_mem[22205] = 0;
disk_mem[22206] = 0;
disk_mem[22207] = 0;
disk_mem[22208] = 0;
disk_mem[22209] = 0;
disk_mem[22210] = 0;
disk_mem[22211] = 0;
disk_mem[22212] = 0;
disk_mem[22213] = 0;
disk_mem[22214] = 0;
disk_mem[22215] = 0;
disk_mem[22216] = 0;
disk_mem[22217] = 0;
disk_mem[22218] = 0;
disk_mem[22219] = 0;
disk_mem[22220] = 0;
disk_mem[22221] = 0;
disk_mem[22222] = 0;
disk_mem[22223] = 0;
disk_mem[22224] = 0;
disk_mem[22225] = 0;
disk_mem[22226] = 0;
disk_mem[22227] = 0;
disk_mem[22228] = 0;
disk_mem[22229] = 0;
disk_mem[22230] = 0;
disk_mem[22231] = 0;
disk_mem[22232] = 0;
disk_mem[22233] = 0;
disk_mem[22234] = 0;
disk_mem[22235] = 0;
disk_mem[22236] = 0;
disk_mem[22237] = 0;
disk_mem[22238] = 0;
disk_mem[22239] = 0;
disk_mem[22240] = 0;
disk_mem[22241] = 0;
disk_mem[22242] = 0;
disk_mem[22243] = 0;
disk_mem[22244] = 0;
disk_mem[22245] = 0;
disk_mem[22246] = 0;
disk_mem[22247] = 0;
disk_mem[22248] = 0;
disk_mem[22249] = 0;
disk_mem[22250] = 0;
disk_mem[22251] = 0;
disk_mem[22252] = 0;
disk_mem[22253] = 0;
disk_mem[22254] = 0;
disk_mem[22255] = 0;
disk_mem[22256] = 0;
disk_mem[22257] = 0;
disk_mem[22258] = 0;
disk_mem[22259] = 0;
disk_mem[22260] = 0;
disk_mem[22261] = 0;
disk_mem[22262] = 0;
disk_mem[22263] = 0;
disk_mem[22264] = 0;
disk_mem[22265] = 0;
disk_mem[22266] = 0;
disk_mem[22267] = 0;
disk_mem[22268] = 0;
disk_mem[22269] = 0;
disk_mem[22270] = 0;
disk_mem[22271] = 0;
disk_mem[22272] = 0;
disk_mem[22273] = 0;
disk_mem[22274] = 0;
disk_mem[22275] = 0;
disk_mem[22276] = 0;
disk_mem[22277] = 0;
disk_mem[22278] = 0;
disk_mem[22279] = 0;
disk_mem[22280] = 0;
disk_mem[22281] = 0;
disk_mem[22282] = 0;
disk_mem[22283] = 0;
disk_mem[22284] = 0;
disk_mem[22285] = 0;
disk_mem[22286] = 0;
disk_mem[22287] = 0;
disk_mem[22288] = 0;
disk_mem[22289] = 0;
disk_mem[22290] = 0;
disk_mem[22291] = 0;
disk_mem[22292] = 0;
disk_mem[22293] = 0;
disk_mem[22294] = 0;
disk_mem[22295] = 0;
disk_mem[22296] = 0;
disk_mem[22297] = 0;
disk_mem[22298] = 0;
disk_mem[22299] = 0;
disk_mem[22300] = 0;
disk_mem[22301] = 0;
disk_mem[22302] = 0;
disk_mem[22303] = 0;
disk_mem[22304] = 0;
disk_mem[22305] = 0;
disk_mem[22306] = 0;
disk_mem[22307] = 0;
disk_mem[22308] = 0;
disk_mem[22309] = 0;
disk_mem[22310] = 0;
disk_mem[22311] = 0;
disk_mem[22312] = 0;
disk_mem[22313] = 0;
disk_mem[22314] = 0;
disk_mem[22315] = 0;
disk_mem[22316] = 0;
disk_mem[22317] = 0;
disk_mem[22318] = 0;
disk_mem[22319] = 0;
disk_mem[22320] = 0;
disk_mem[22321] = 0;
disk_mem[22322] = 0;
disk_mem[22323] = 0;
disk_mem[22324] = 0;
disk_mem[22325] = 0;
disk_mem[22326] = 0;
disk_mem[22327] = 0;
disk_mem[22328] = 0;
disk_mem[22329] = 0;
disk_mem[22330] = 0;
disk_mem[22331] = 0;
disk_mem[22332] = 0;
disk_mem[22333] = 0;
disk_mem[22334] = 0;
disk_mem[22335] = 0;
disk_mem[22336] = 0;
disk_mem[22337] = 0;
disk_mem[22338] = 0;
disk_mem[22339] = 0;
disk_mem[22340] = 0;
disk_mem[22341] = 0;
disk_mem[22342] = 0;
disk_mem[22343] = 0;
disk_mem[22344] = 0;
disk_mem[22345] = 0;
disk_mem[22346] = 0;
disk_mem[22347] = 0;
disk_mem[22348] = 0;
disk_mem[22349] = 0;
disk_mem[22350] = 0;
disk_mem[22351] = 0;
disk_mem[22352] = 0;
disk_mem[22353] = 0;
disk_mem[22354] = 0;
disk_mem[22355] = 0;
disk_mem[22356] = 0;
disk_mem[22357] = 0;
disk_mem[22358] = 0;
disk_mem[22359] = 0;
disk_mem[22360] = 0;
disk_mem[22361] = 0;
disk_mem[22362] = 0;
disk_mem[22363] = 0;
disk_mem[22364] = 0;
disk_mem[22365] = 0;
disk_mem[22366] = 0;
disk_mem[22367] = 0;
disk_mem[22368] = 0;
disk_mem[22369] = 0;
disk_mem[22370] = 0;
disk_mem[22371] = 0;
disk_mem[22372] = 0;
disk_mem[22373] = 0;
disk_mem[22374] = 0;
disk_mem[22375] = 0;
disk_mem[22376] = 0;
disk_mem[22377] = 0;
disk_mem[22378] = 0;
disk_mem[22379] = 0;
disk_mem[22380] = 0;
disk_mem[22381] = 0;
disk_mem[22382] = 0;
disk_mem[22383] = 0;
disk_mem[22384] = 0;
disk_mem[22385] = 0;
disk_mem[22386] = 0;
disk_mem[22387] = 0;
disk_mem[22388] = 0;
disk_mem[22389] = 0;
disk_mem[22390] = 0;
disk_mem[22391] = 0;
disk_mem[22392] = 0;
disk_mem[22393] = 0;
disk_mem[22394] = 0;
disk_mem[22395] = 0;
disk_mem[22396] = 0;
disk_mem[22397] = 0;
disk_mem[22398] = 0;
disk_mem[22399] = 0;
disk_mem[22400] = 0;
disk_mem[22401] = 0;
disk_mem[22402] = 0;
disk_mem[22403] = 0;
disk_mem[22404] = 0;
disk_mem[22405] = 0;
disk_mem[22406] = 0;
disk_mem[22407] = 0;
disk_mem[22408] = 0;
disk_mem[22409] = 0;
disk_mem[22410] = 0;
disk_mem[22411] = 0;
disk_mem[22412] = 0;
disk_mem[22413] = 0;
disk_mem[22414] = 0;
disk_mem[22415] = 0;
disk_mem[22416] = 0;
disk_mem[22417] = 0;
disk_mem[22418] = 0;
disk_mem[22419] = 0;
disk_mem[22420] = 0;
disk_mem[22421] = 0;
disk_mem[22422] = 0;
disk_mem[22423] = 0;
disk_mem[22424] = 0;
disk_mem[22425] = 0;
disk_mem[22426] = 0;
disk_mem[22427] = 0;
disk_mem[22428] = 0;
disk_mem[22429] = 0;
disk_mem[22430] = 0;
disk_mem[22431] = 0;
disk_mem[22432] = 0;
disk_mem[22433] = 0;
disk_mem[22434] = 0;
disk_mem[22435] = 0;
disk_mem[22436] = 0;
disk_mem[22437] = 0;
disk_mem[22438] = 0;
disk_mem[22439] = 0;
disk_mem[22440] = 0;
disk_mem[22441] = 0;
disk_mem[22442] = 0;
disk_mem[22443] = 0;
disk_mem[22444] = 0;
disk_mem[22445] = 0;
disk_mem[22446] = 0;
disk_mem[22447] = 0;
disk_mem[22448] = 0;
disk_mem[22449] = 0;
disk_mem[22450] = 0;
disk_mem[22451] = 0;
disk_mem[22452] = 0;
disk_mem[22453] = 0;
disk_mem[22454] = 0;
disk_mem[22455] = 0;
disk_mem[22456] = 0;
disk_mem[22457] = 0;
disk_mem[22458] = 0;
disk_mem[22459] = 0;
disk_mem[22460] = 0;
disk_mem[22461] = 0;
disk_mem[22462] = 0;
disk_mem[22463] = 0;
disk_mem[22464] = 0;
disk_mem[22465] = 0;
disk_mem[22466] = 0;
disk_mem[22467] = 0;
disk_mem[22468] = 0;
disk_mem[22469] = 0;
disk_mem[22470] = 0;
disk_mem[22471] = 0;
disk_mem[22472] = 0;
disk_mem[22473] = 0;
disk_mem[22474] = 0;
disk_mem[22475] = 0;
disk_mem[22476] = 0;
disk_mem[22477] = 0;
disk_mem[22478] = 0;
disk_mem[22479] = 0;
disk_mem[22480] = 0;
disk_mem[22481] = 0;
disk_mem[22482] = 0;
disk_mem[22483] = 0;
disk_mem[22484] = 0;
disk_mem[22485] = 0;
disk_mem[22486] = 0;
disk_mem[22487] = 0;
disk_mem[22488] = 0;
disk_mem[22489] = 0;
disk_mem[22490] = 0;
disk_mem[22491] = 0;
disk_mem[22492] = 0;
disk_mem[22493] = 0;
disk_mem[22494] = 0;
disk_mem[22495] = 0;
disk_mem[22496] = 0;
disk_mem[22497] = 0;
disk_mem[22498] = 0;
disk_mem[22499] = 0;
disk_mem[22500] = 0;
disk_mem[22501] = 0;
disk_mem[22502] = 0;
disk_mem[22503] = 0;
disk_mem[22504] = 0;
disk_mem[22505] = 0;
disk_mem[22506] = 0;
disk_mem[22507] = 0;
disk_mem[22508] = 0;
disk_mem[22509] = 0;
disk_mem[22510] = 0;
disk_mem[22511] = 0;
disk_mem[22512] = 0;
disk_mem[22513] = 0;
disk_mem[22514] = 0;
disk_mem[22515] = 0;
disk_mem[22516] = 0;
disk_mem[22517] = 0;
disk_mem[22518] = 0;
disk_mem[22519] = 0;
disk_mem[22520] = 0;
disk_mem[22521] = 0;
disk_mem[22522] = 0;
disk_mem[22523] = 0;
disk_mem[22524] = 0;
disk_mem[22525] = 0;
disk_mem[22526] = 0;
disk_mem[22527] = 0;
disk_mem[22528] = 'h48;
disk_mem[22529] = 'h65;
disk_mem[22530] = 'h6C;
disk_mem[22531] = 'h6C;
disk_mem[22532] = 'h6F;
disk_mem[22533] = 'h20;
disk_mem[22534] = 'h77;
disk_mem[22535] = 'h6F;
disk_mem[22536] = 'h72;
disk_mem[22537] = 'h6C;
disk_mem[22538] = 'h64;
disk_mem[22539] = 'h21;
disk_mem[22540] = 'h0D;
disk_mem[22541] = 'h0A;
disk_mem[22542] = 'h41;
disk_mem[22543] = 'h20;
disk_mem[22544] = 'h32;
disk_mem[22545] = 'h34;
disk_mem[22546] = 'h6B;
disk_mem[22547] = 'h42;
disk_mem[22548] = 'h20;
disk_mem[22549] = 'h64;
disk_mem[22550] = 'h69;
disk_mem[22551] = 'h73;
disk_mem[22552] = 'h6B;
disk_mem[22553] = 'h20;
disk_mem[22554] = 'h70;
disk_mem[22555] = 'h61;
disk_mem[22556] = 'h72;
disk_mem[22557] = 'h74;
disk_mem[22558] = 'h69;
disk_mem[22559] = 'h74;
disk_mem[22560] = 'h69;
disk_mem[22561] = 'h6F;
disk_mem[22562] = 'h6E;
disk_mem[22563] = 'h2E;
disk_mem[22564] = 'h0D;
disk_mem[22565] = 'h0A;
disk_mem[22566] = 0;
disk_mem[22567] = 0;
disk_mem[22568] = 0;
disk_mem[22569] = 0;
disk_mem[22570] = 0;
disk_mem[22571] = 0;
disk_mem[22572] = 0;
disk_mem[22573] = 0;
disk_mem[22574] = 0;
disk_mem[22575] = 0;
disk_mem[22576] = 0;
disk_mem[22577] = 0;
disk_mem[22578] = 0;
disk_mem[22579] = 0;
disk_mem[22580] = 0;
disk_mem[22581] = 0;
disk_mem[22582] = 0;
disk_mem[22583] = 0;
disk_mem[22584] = 0;
disk_mem[22585] = 0;
disk_mem[22586] = 0;
disk_mem[22587] = 0;
disk_mem[22588] = 0;
disk_mem[22589] = 0;
disk_mem[22590] = 0;
disk_mem[22591] = 0;
disk_mem[22592] = 0;
disk_mem[22593] = 0;
disk_mem[22594] = 0;
disk_mem[22595] = 0;
disk_mem[22596] = 0;
disk_mem[22597] = 0;
disk_mem[22598] = 0;
disk_mem[22599] = 0;
disk_mem[22600] = 0;
disk_mem[22601] = 0;
disk_mem[22602] = 0;
disk_mem[22603] = 0;
disk_mem[22604] = 0;
disk_mem[22605] = 0;
disk_mem[22606] = 0;
disk_mem[22607] = 0;
disk_mem[22608] = 0;
disk_mem[22609] = 0;
disk_mem[22610] = 0;
disk_mem[22611] = 0;
disk_mem[22612] = 0;
disk_mem[22613] = 0;
disk_mem[22614] = 0;
disk_mem[22615] = 0;
disk_mem[22616] = 0;
disk_mem[22617] = 0;
disk_mem[22618] = 0;
disk_mem[22619] = 0;
disk_mem[22620] = 0;
disk_mem[22621] = 0;
disk_mem[22622] = 0;
disk_mem[22623] = 0;
disk_mem[22624] = 0;
disk_mem[22625] = 0;
disk_mem[22626] = 0;
disk_mem[22627] = 0;
disk_mem[22628] = 0;
disk_mem[22629] = 0;
disk_mem[22630] = 0;
disk_mem[22631] = 0;
disk_mem[22632] = 0;
disk_mem[22633] = 0;
disk_mem[22634] = 0;
disk_mem[22635] = 0;
disk_mem[22636] = 0;
disk_mem[22637] = 0;
disk_mem[22638] = 0;
disk_mem[22639] = 0;
disk_mem[22640] = 0;
disk_mem[22641] = 0;
disk_mem[22642] = 0;
disk_mem[22643] = 0;
disk_mem[22644] = 0;
disk_mem[22645] = 0;
disk_mem[22646] = 0;
disk_mem[22647] = 0;
disk_mem[22648] = 0;
disk_mem[22649] = 0;
disk_mem[22650] = 0;
disk_mem[22651] = 0;
disk_mem[22652] = 0;
disk_mem[22653] = 0;
disk_mem[22654] = 0;
disk_mem[22655] = 0;
disk_mem[22656] = 0;
disk_mem[22657] = 0;
disk_mem[22658] = 0;
disk_mem[22659] = 0;
disk_mem[22660] = 0;
disk_mem[22661] = 0;
disk_mem[22662] = 0;
disk_mem[22663] = 0;
disk_mem[22664] = 0;
disk_mem[22665] = 0;
disk_mem[22666] = 0;
disk_mem[22667] = 0;
disk_mem[22668] = 0;
disk_mem[22669] = 0;
disk_mem[22670] = 0;
disk_mem[22671] = 0;
disk_mem[22672] = 0;
disk_mem[22673] = 0;
disk_mem[22674] = 0;
disk_mem[22675] = 0;
disk_mem[22676] = 0;
disk_mem[22677] = 0;
disk_mem[22678] = 0;
disk_mem[22679] = 0;
disk_mem[22680] = 0;
disk_mem[22681] = 0;
disk_mem[22682] = 0;
disk_mem[22683] = 0;
disk_mem[22684] = 0;
disk_mem[22685] = 0;
disk_mem[22686] = 0;
disk_mem[22687] = 0;
disk_mem[22688] = 0;
disk_mem[22689] = 0;
disk_mem[22690] = 0;
disk_mem[22691] = 0;
disk_mem[22692] = 0;
disk_mem[22693] = 0;
disk_mem[22694] = 0;
disk_mem[22695] = 0;
disk_mem[22696] = 0;
disk_mem[22697] = 0;
disk_mem[22698] = 0;
disk_mem[22699] = 0;
disk_mem[22700] = 0;
disk_mem[22701] = 0;
disk_mem[22702] = 0;
disk_mem[22703] = 0;
disk_mem[22704] = 0;
disk_mem[22705] = 0;
disk_mem[22706] = 0;
disk_mem[22707] = 0;
disk_mem[22708] = 0;
disk_mem[22709] = 0;
disk_mem[22710] = 0;
disk_mem[22711] = 0;
disk_mem[22712] = 0;
disk_mem[22713] = 0;
disk_mem[22714] = 0;
disk_mem[22715] = 0;
disk_mem[22716] = 0;
disk_mem[22717] = 0;
disk_mem[22718] = 0;
disk_mem[22719] = 0;
disk_mem[22720] = 0;
disk_mem[22721] = 0;
disk_mem[22722] = 0;
disk_mem[22723] = 0;
disk_mem[22724] = 0;
disk_mem[22725] = 0;
disk_mem[22726] = 0;
disk_mem[22727] = 0;
disk_mem[22728] = 0;
disk_mem[22729] = 0;
disk_mem[22730] = 0;
disk_mem[22731] = 0;
disk_mem[22732] = 0;
disk_mem[22733] = 0;
disk_mem[22734] = 0;
disk_mem[22735] = 0;
disk_mem[22736] = 0;
disk_mem[22737] = 0;
disk_mem[22738] = 0;
disk_mem[22739] = 0;
disk_mem[22740] = 0;
disk_mem[22741] = 0;
disk_mem[22742] = 0;
disk_mem[22743] = 0;
disk_mem[22744] = 0;
disk_mem[22745] = 0;
disk_mem[22746] = 0;
disk_mem[22747] = 0;
disk_mem[22748] = 0;
disk_mem[22749] = 0;
disk_mem[22750] = 0;
disk_mem[22751] = 0;
disk_mem[22752] = 0;
disk_mem[22753] = 0;
disk_mem[22754] = 0;
disk_mem[22755] = 0;
disk_mem[22756] = 0;
disk_mem[22757] = 0;
disk_mem[22758] = 0;
disk_mem[22759] = 0;
disk_mem[22760] = 0;
disk_mem[22761] = 0;
disk_mem[22762] = 0;
disk_mem[22763] = 0;
disk_mem[22764] = 0;
disk_mem[22765] = 0;
disk_mem[22766] = 0;
disk_mem[22767] = 0;
disk_mem[22768] = 0;
disk_mem[22769] = 0;
disk_mem[22770] = 0;
disk_mem[22771] = 0;
disk_mem[22772] = 0;
disk_mem[22773] = 0;
disk_mem[22774] = 0;
disk_mem[22775] = 0;
disk_mem[22776] = 0;
disk_mem[22777] = 0;
disk_mem[22778] = 0;
disk_mem[22779] = 0;
disk_mem[22780] = 0;
disk_mem[22781] = 0;
disk_mem[22782] = 0;
disk_mem[22783] = 0;
disk_mem[22784] = 0;
disk_mem[22785] = 0;
disk_mem[22786] = 0;
disk_mem[22787] = 0;
disk_mem[22788] = 0;
disk_mem[22789] = 0;
disk_mem[22790] = 0;
disk_mem[22791] = 0;
disk_mem[22792] = 0;
disk_mem[22793] = 0;
disk_mem[22794] = 0;
disk_mem[22795] = 0;
disk_mem[22796] = 0;
disk_mem[22797] = 0;
disk_mem[22798] = 0;
disk_mem[22799] = 0;
disk_mem[22800] = 0;
disk_mem[22801] = 0;
disk_mem[22802] = 0;
disk_mem[22803] = 0;
disk_mem[22804] = 0;
disk_mem[22805] = 0;
disk_mem[22806] = 0;
disk_mem[22807] = 0;
disk_mem[22808] = 0;
disk_mem[22809] = 0;
disk_mem[22810] = 0;
disk_mem[22811] = 0;
disk_mem[22812] = 0;
disk_mem[22813] = 0;
disk_mem[22814] = 0;
disk_mem[22815] = 0;
disk_mem[22816] = 0;
disk_mem[22817] = 0;
disk_mem[22818] = 0;
disk_mem[22819] = 0;
disk_mem[22820] = 0;
disk_mem[22821] = 0;
disk_mem[22822] = 0;
disk_mem[22823] = 0;
disk_mem[22824] = 0;
disk_mem[22825] = 0;
disk_mem[22826] = 0;
disk_mem[22827] = 0;
disk_mem[22828] = 0;
disk_mem[22829] = 0;
disk_mem[22830] = 0;
disk_mem[22831] = 0;
disk_mem[22832] = 0;
disk_mem[22833] = 0;
disk_mem[22834] = 0;
disk_mem[22835] = 0;
disk_mem[22836] = 0;
disk_mem[22837] = 0;
disk_mem[22838] = 0;
disk_mem[22839] = 0;
disk_mem[22840] = 0;
disk_mem[22841] = 0;
disk_mem[22842] = 0;
disk_mem[22843] = 0;
disk_mem[22844] = 0;
disk_mem[22845] = 0;
disk_mem[22846] = 0;
disk_mem[22847] = 0;
disk_mem[22848] = 0;
disk_mem[22849] = 0;
disk_mem[22850] = 0;
disk_mem[22851] = 0;
disk_mem[22852] = 0;
disk_mem[22853] = 0;
disk_mem[22854] = 0;
disk_mem[22855] = 0;
disk_mem[22856] = 0;
disk_mem[22857] = 0;
disk_mem[22858] = 0;
disk_mem[22859] = 0;
disk_mem[22860] = 0;
disk_mem[22861] = 0;
disk_mem[22862] = 0;
disk_mem[22863] = 0;
disk_mem[22864] = 0;
disk_mem[22865] = 0;
disk_mem[22866] = 0;
disk_mem[22867] = 0;
disk_mem[22868] = 0;
disk_mem[22869] = 0;
disk_mem[22870] = 0;
disk_mem[22871] = 0;
disk_mem[22872] = 0;
disk_mem[22873] = 0;
disk_mem[22874] = 0;
disk_mem[22875] = 0;
disk_mem[22876] = 0;
disk_mem[22877] = 0;
disk_mem[22878] = 0;
disk_mem[22879] = 0;
disk_mem[22880] = 0;
disk_mem[22881] = 0;
disk_mem[22882] = 0;
disk_mem[22883] = 0;
disk_mem[22884] = 0;
disk_mem[22885] = 0;
disk_mem[22886] = 0;
disk_mem[22887] = 0;
disk_mem[22888] = 0;
disk_mem[22889] = 0;
disk_mem[22890] = 0;
disk_mem[22891] = 0;
disk_mem[22892] = 0;
disk_mem[22893] = 0;
disk_mem[22894] = 0;
disk_mem[22895] = 0;
disk_mem[22896] = 0;
disk_mem[22897] = 0;
disk_mem[22898] = 0;
disk_mem[22899] = 0;
disk_mem[22900] = 0;
disk_mem[22901] = 0;
disk_mem[22902] = 0;
disk_mem[22903] = 0;
disk_mem[22904] = 0;
disk_mem[22905] = 0;
disk_mem[22906] = 0;
disk_mem[22907] = 0;
disk_mem[22908] = 0;
disk_mem[22909] = 0;
disk_mem[22910] = 0;
disk_mem[22911] = 0;
disk_mem[22912] = 0;
disk_mem[22913] = 0;
disk_mem[22914] = 0;
disk_mem[22915] = 0;
disk_mem[22916] = 0;
disk_mem[22917] = 0;
disk_mem[22918] = 0;
disk_mem[22919] = 0;
disk_mem[22920] = 0;
disk_mem[22921] = 0;
disk_mem[22922] = 0;
disk_mem[22923] = 0;
disk_mem[22924] = 0;
disk_mem[22925] = 0;
disk_mem[22926] = 0;
disk_mem[22927] = 0;
disk_mem[22928] = 0;
disk_mem[22929] = 0;
disk_mem[22930] = 0;
disk_mem[22931] = 0;
disk_mem[22932] = 0;
disk_mem[22933] = 0;
disk_mem[22934] = 0;
disk_mem[22935] = 0;
disk_mem[22936] = 0;
disk_mem[22937] = 0;
disk_mem[22938] = 0;
disk_mem[22939] = 0;
disk_mem[22940] = 0;
disk_mem[22941] = 0;
disk_mem[22942] = 0;
disk_mem[22943] = 0;
disk_mem[22944] = 0;
disk_mem[22945] = 0;
disk_mem[22946] = 0;
disk_mem[22947] = 0;
disk_mem[22948] = 0;
disk_mem[22949] = 0;
disk_mem[22950] = 0;
disk_mem[22951] = 0;
disk_mem[22952] = 0;
disk_mem[22953] = 0;
disk_mem[22954] = 0;
disk_mem[22955] = 0;
disk_mem[22956] = 0;
disk_mem[22957] = 0;
disk_mem[22958] = 0;
disk_mem[22959] = 0;
disk_mem[22960] = 0;
disk_mem[22961] = 0;
disk_mem[22962] = 0;
disk_mem[22963] = 0;
disk_mem[22964] = 0;
disk_mem[22965] = 0;
disk_mem[22966] = 0;
disk_mem[22967] = 0;
disk_mem[22968] = 0;
disk_mem[22969] = 0;
disk_mem[22970] = 0;
disk_mem[22971] = 0;
disk_mem[22972] = 0;
disk_mem[22973] = 0;
disk_mem[22974] = 0;
disk_mem[22975] = 0;
disk_mem[22976] = 0;
disk_mem[22977] = 0;
disk_mem[22978] = 0;
disk_mem[22979] = 0;
disk_mem[22980] = 0;
disk_mem[22981] = 0;
disk_mem[22982] = 0;
disk_mem[22983] = 0;
disk_mem[22984] = 0;
disk_mem[22985] = 0;
disk_mem[22986] = 0;
disk_mem[22987] = 0;
disk_mem[22988] = 0;
disk_mem[22989] = 0;
disk_mem[22990] = 0;
disk_mem[22991] = 0;
disk_mem[22992] = 0;
disk_mem[22993] = 0;
disk_mem[22994] = 0;
disk_mem[22995] = 0;
disk_mem[22996] = 0;
disk_mem[22997] = 0;
disk_mem[22998] = 0;
disk_mem[22999] = 0;
disk_mem[23000] = 0;
disk_mem[23001] = 0;
disk_mem[23002] = 0;
disk_mem[23003] = 0;
disk_mem[23004] = 0;
disk_mem[23005] = 0;
disk_mem[23006] = 0;
disk_mem[23007] = 0;
disk_mem[23008] = 0;
disk_mem[23009] = 0;
disk_mem[23010] = 0;
disk_mem[23011] = 0;
disk_mem[23012] = 0;
disk_mem[23013] = 0;
disk_mem[23014] = 0;
disk_mem[23015] = 0;
disk_mem[23016] = 0;
disk_mem[23017] = 0;
disk_mem[23018] = 0;
disk_mem[23019] = 0;
disk_mem[23020] = 0;
disk_mem[23021] = 0;
disk_mem[23022] = 0;
disk_mem[23023] = 0;
disk_mem[23024] = 0;
disk_mem[23025] = 0;
disk_mem[23026] = 0;
disk_mem[23027] = 0;
disk_mem[23028] = 0;
disk_mem[23029] = 0;
disk_mem[23030] = 0;
disk_mem[23031] = 0;
disk_mem[23032] = 0;
disk_mem[23033] = 0;
disk_mem[23034] = 0;
disk_mem[23035] = 0;
disk_mem[23036] = 0;
disk_mem[23037] = 0;
disk_mem[23038] = 0;
disk_mem[23039] = 0;
disk_mem[23040] = 0;
disk_mem[23041] = 0;
disk_mem[23042] = 0;
disk_mem[23043] = 0;
disk_mem[23044] = 0;
disk_mem[23045] = 0;
disk_mem[23046] = 0;
disk_mem[23047] = 0;
disk_mem[23048] = 0;
disk_mem[23049] = 0;
disk_mem[23050] = 0;
disk_mem[23051] = 0;
disk_mem[23052] = 0;
disk_mem[23053] = 0;
disk_mem[23054] = 0;
disk_mem[23055] = 0;
disk_mem[23056] = 0;
disk_mem[23057] = 0;
disk_mem[23058] = 0;
disk_mem[23059] = 0;
disk_mem[23060] = 0;
disk_mem[23061] = 0;
disk_mem[23062] = 0;
disk_mem[23063] = 0;
disk_mem[23064] = 0;
disk_mem[23065] = 0;
disk_mem[23066] = 0;
disk_mem[23067] = 0;
disk_mem[23068] = 0;
disk_mem[23069] = 0;
disk_mem[23070] = 0;
disk_mem[23071] = 0;
disk_mem[23072] = 0;
disk_mem[23073] = 0;
disk_mem[23074] = 0;
disk_mem[23075] = 0;
disk_mem[23076] = 0;
disk_mem[23077] = 0;
disk_mem[23078] = 0;
disk_mem[23079] = 0;
disk_mem[23080] = 0;
disk_mem[23081] = 0;
disk_mem[23082] = 0;
disk_mem[23083] = 0;
disk_mem[23084] = 0;
disk_mem[23085] = 0;
disk_mem[23086] = 0;
disk_mem[23087] = 0;
disk_mem[23088] = 0;
disk_mem[23089] = 0;
disk_mem[23090] = 0;
disk_mem[23091] = 0;
disk_mem[23092] = 0;
disk_mem[23093] = 0;
disk_mem[23094] = 0;
disk_mem[23095] = 0;
disk_mem[23096] = 0;
disk_mem[23097] = 0;
disk_mem[23098] = 0;
disk_mem[23099] = 0;
disk_mem[23100] = 0;
disk_mem[23101] = 0;
disk_mem[23102] = 0;
disk_mem[23103] = 0;
disk_mem[23104] = 0;
disk_mem[23105] = 0;
disk_mem[23106] = 0;
disk_mem[23107] = 0;
disk_mem[23108] = 0;
disk_mem[23109] = 0;
disk_mem[23110] = 0;
disk_mem[23111] = 0;
disk_mem[23112] = 0;
disk_mem[23113] = 0;
disk_mem[23114] = 0;
disk_mem[23115] = 0;
disk_mem[23116] = 0;
disk_mem[23117] = 0;
disk_mem[23118] = 0;
disk_mem[23119] = 0;
disk_mem[23120] = 0;
disk_mem[23121] = 0;
disk_mem[23122] = 0;
disk_mem[23123] = 0;
disk_mem[23124] = 0;
disk_mem[23125] = 0;
disk_mem[23126] = 0;
disk_mem[23127] = 0;
disk_mem[23128] = 0;
disk_mem[23129] = 0;
disk_mem[23130] = 0;
disk_mem[23131] = 0;
disk_mem[23132] = 0;
disk_mem[23133] = 0;
disk_mem[23134] = 0;
disk_mem[23135] = 0;
disk_mem[23136] = 0;
disk_mem[23137] = 0;
disk_mem[23138] = 0;
disk_mem[23139] = 0;
disk_mem[23140] = 0;
disk_mem[23141] = 0;
disk_mem[23142] = 0;
disk_mem[23143] = 0;
disk_mem[23144] = 0;
disk_mem[23145] = 0;
disk_mem[23146] = 0;
disk_mem[23147] = 0;
disk_mem[23148] = 0;
disk_mem[23149] = 0;
disk_mem[23150] = 0;
disk_mem[23151] = 0;
disk_mem[23152] = 0;
disk_mem[23153] = 0;
disk_mem[23154] = 0;
disk_mem[23155] = 0;
disk_mem[23156] = 0;
disk_mem[23157] = 0;
disk_mem[23158] = 0;
disk_mem[23159] = 0;
disk_mem[23160] = 0;
disk_mem[23161] = 0;
disk_mem[23162] = 0;
disk_mem[23163] = 0;
disk_mem[23164] = 0;
disk_mem[23165] = 0;
disk_mem[23166] = 0;
disk_mem[23167] = 0;
disk_mem[23168] = 0;
disk_mem[23169] = 0;
disk_mem[23170] = 0;
disk_mem[23171] = 0;
disk_mem[23172] = 0;
disk_mem[23173] = 0;
disk_mem[23174] = 0;
disk_mem[23175] = 0;
disk_mem[23176] = 0;
disk_mem[23177] = 0;
disk_mem[23178] = 0;
disk_mem[23179] = 0;
disk_mem[23180] = 0;
disk_mem[23181] = 0;
disk_mem[23182] = 0;
disk_mem[23183] = 0;
disk_mem[23184] = 0;
disk_mem[23185] = 0;
disk_mem[23186] = 0;
disk_mem[23187] = 0;
disk_mem[23188] = 0;
disk_mem[23189] = 0;
disk_mem[23190] = 0;
disk_mem[23191] = 0;
disk_mem[23192] = 0;
disk_mem[23193] = 0;
disk_mem[23194] = 0;
disk_mem[23195] = 0;
disk_mem[23196] = 0;
disk_mem[23197] = 0;
disk_mem[23198] = 0;
disk_mem[23199] = 0;
disk_mem[23200] = 0;
disk_mem[23201] = 0;
disk_mem[23202] = 0;
disk_mem[23203] = 0;
disk_mem[23204] = 0;
disk_mem[23205] = 0;
disk_mem[23206] = 0;
disk_mem[23207] = 0;
disk_mem[23208] = 0;
disk_mem[23209] = 0;
disk_mem[23210] = 0;
disk_mem[23211] = 0;
disk_mem[23212] = 0;
disk_mem[23213] = 0;
disk_mem[23214] = 0;
disk_mem[23215] = 0;
disk_mem[23216] = 0;
disk_mem[23217] = 0;
disk_mem[23218] = 0;
disk_mem[23219] = 0;
disk_mem[23220] = 0;
disk_mem[23221] = 0;
disk_mem[23222] = 0;
disk_mem[23223] = 0;
disk_mem[23224] = 0;
disk_mem[23225] = 0;
disk_mem[23226] = 0;
disk_mem[23227] = 0;
disk_mem[23228] = 0;
disk_mem[23229] = 0;
disk_mem[23230] = 0;
disk_mem[23231] = 0;
disk_mem[23232] = 0;
disk_mem[23233] = 0;
disk_mem[23234] = 0;
disk_mem[23235] = 0;
disk_mem[23236] = 0;
disk_mem[23237] = 0;
disk_mem[23238] = 0;
disk_mem[23239] = 0;
disk_mem[23240] = 0;
disk_mem[23241] = 0;
disk_mem[23242] = 0;
disk_mem[23243] = 0;
disk_mem[23244] = 0;
disk_mem[23245] = 0;
disk_mem[23246] = 0;
disk_mem[23247] = 0;
disk_mem[23248] = 0;
disk_mem[23249] = 0;
disk_mem[23250] = 0;
disk_mem[23251] = 0;
disk_mem[23252] = 0;
disk_mem[23253] = 0;
disk_mem[23254] = 0;
disk_mem[23255] = 0;
disk_mem[23256] = 0;
disk_mem[23257] = 0;
disk_mem[23258] = 0;
disk_mem[23259] = 0;
disk_mem[23260] = 0;
disk_mem[23261] = 0;
disk_mem[23262] = 0;
disk_mem[23263] = 0;
disk_mem[23264] = 0;
disk_mem[23265] = 0;
disk_mem[23266] = 0;
disk_mem[23267] = 0;
disk_mem[23268] = 0;
disk_mem[23269] = 0;
disk_mem[23270] = 0;
disk_mem[23271] = 0;
disk_mem[23272] = 0;
disk_mem[23273] = 0;
disk_mem[23274] = 0;
disk_mem[23275] = 0;
disk_mem[23276] = 0;
disk_mem[23277] = 0;
disk_mem[23278] = 0;
disk_mem[23279] = 0;
disk_mem[23280] = 0;
disk_mem[23281] = 0;
disk_mem[23282] = 0;
disk_mem[23283] = 0;
disk_mem[23284] = 0;
disk_mem[23285] = 0;
disk_mem[23286] = 0;
disk_mem[23287] = 0;
disk_mem[23288] = 0;
disk_mem[23289] = 0;
disk_mem[23290] = 0;
disk_mem[23291] = 0;
disk_mem[23292] = 0;
disk_mem[23293] = 0;
disk_mem[23294] = 0;
disk_mem[23295] = 0;
disk_mem[23296] = 0;
disk_mem[23297] = 0;
disk_mem[23298] = 0;
disk_mem[23299] = 0;
disk_mem[23300] = 0;
disk_mem[23301] = 0;
disk_mem[23302] = 0;
disk_mem[23303] = 0;
disk_mem[23304] = 0;
disk_mem[23305] = 0;
disk_mem[23306] = 0;
disk_mem[23307] = 0;
disk_mem[23308] = 0;
disk_mem[23309] = 0;
disk_mem[23310] = 0;
disk_mem[23311] = 0;
disk_mem[23312] = 0;
disk_mem[23313] = 0;
disk_mem[23314] = 0;
disk_mem[23315] = 0;
disk_mem[23316] = 0;
disk_mem[23317] = 0;
disk_mem[23318] = 0;
disk_mem[23319] = 0;
disk_mem[23320] = 0;
disk_mem[23321] = 0;
disk_mem[23322] = 0;
disk_mem[23323] = 0;
disk_mem[23324] = 0;
disk_mem[23325] = 0;
disk_mem[23326] = 0;
disk_mem[23327] = 0;
disk_mem[23328] = 0;
disk_mem[23329] = 0;
disk_mem[23330] = 0;
disk_mem[23331] = 0;
disk_mem[23332] = 0;
disk_mem[23333] = 0;
disk_mem[23334] = 0;
disk_mem[23335] = 0;
disk_mem[23336] = 0;
disk_mem[23337] = 0;
disk_mem[23338] = 0;
disk_mem[23339] = 0;
disk_mem[23340] = 0;
disk_mem[23341] = 0;
disk_mem[23342] = 0;
disk_mem[23343] = 0;
disk_mem[23344] = 0;
disk_mem[23345] = 0;
disk_mem[23346] = 0;
disk_mem[23347] = 0;
disk_mem[23348] = 0;
disk_mem[23349] = 0;
disk_mem[23350] = 0;
disk_mem[23351] = 0;
disk_mem[23352] = 0;
disk_mem[23353] = 0;
disk_mem[23354] = 0;
disk_mem[23355] = 0;
disk_mem[23356] = 0;
disk_mem[23357] = 0;
disk_mem[23358] = 0;
disk_mem[23359] = 0;
disk_mem[23360] = 0;
disk_mem[23361] = 0;
disk_mem[23362] = 0;
disk_mem[23363] = 0;
disk_mem[23364] = 0;
disk_mem[23365] = 0;
disk_mem[23366] = 0;
disk_mem[23367] = 0;
disk_mem[23368] = 0;
disk_mem[23369] = 0;
disk_mem[23370] = 0;
disk_mem[23371] = 0;
disk_mem[23372] = 0;
disk_mem[23373] = 0;
disk_mem[23374] = 0;
disk_mem[23375] = 0;
disk_mem[23376] = 0;
disk_mem[23377] = 0;
disk_mem[23378] = 0;
disk_mem[23379] = 0;
disk_mem[23380] = 0;
disk_mem[23381] = 0;
disk_mem[23382] = 0;
disk_mem[23383] = 0;
disk_mem[23384] = 0;
disk_mem[23385] = 0;
disk_mem[23386] = 0;
disk_mem[23387] = 0;
disk_mem[23388] = 0;
disk_mem[23389] = 0;
disk_mem[23390] = 0;
disk_mem[23391] = 0;
disk_mem[23392] = 0;
disk_mem[23393] = 0;
disk_mem[23394] = 0;
disk_mem[23395] = 0;
disk_mem[23396] = 0;
disk_mem[23397] = 0;
disk_mem[23398] = 0;
disk_mem[23399] = 0;
disk_mem[23400] = 0;
disk_mem[23401] = 0;
disk_mem[23402] = 0;
disk_mem[23403] = 0;
disk_mem[23404] = 0;
disk_mem[23405] = 0;
disk_mem[23406] = 0;
disk_mem[23407] = 0;
disk_mem[23408] = 0;
disk_mem[23409] = 0;
disk_mem[23410] = 0;
disk_mem[23411] = 0;
disk_mem[23412] = 0;
disk_mem[23413] = 0;
disk_mem[23414] = 0;
disk_mem[23415] = 0;
disk_mem[23416] = 0;
disk_mem[23417] = 0;
disk_mem[23418] = 0;
disk_mem[23419] = 0;
disk_mem[23420] = 0;
disk_mem[23421] = 0;
disk_mem[23422] = 0;
disk_mem[23423] = 0;
disk_mem[23424] = 0;
disk_mem[23425] = 0;
disk_mem[23426] = 0;
disk_mem[23427] = 0;
disk_mem[23428] = 0;
disk_mem[23429] = 0;
disk_mem[23430] = 0;
disk_mem[23431] = 0;
disk_mem[23432] = 0;
disk_mem[23433] = 0;
disk_mem[23434] = 0;
disk_mem[23435] = 0;
disk_mem[23436] = 0;
disk_mem[23437] = 0;
disk_mem[23438] = 0;
disk_mem[23439] = 0;
disk_mem[23440] = 0;
disk_mem[23441] = 0;
disk_mem[23442] = 0;
disk_mem[23443] = 0;
disk_mem[23444] = 0;
disk_mem[23445] = 0;
disk_mem[23446] = 0;
disk_mem[23447] = 0;
disk_mem[23448] = 0;
disk_mem[23449] = 0;
disk_mem[23450] = 0;
disk_mem[23451] = 0;
disk_mem[23452] = 0;
disk_mem[23453] = 0;
disk_mem[23454] = 0;
disk_mem[23455] = 0;
disk_mem[23456] = 0;
disk_mem[23457] = 0;
disk_mem[23458] = 0;
disk_mem[23459] = 0;
disk_mem[23460] = 0;
disk_mem[23461] = 0;
disk_mem[23462] = 0;
disk_mem[23463] = 0;
disk_mem[23464] = 0;
disk_mem[23465] = 0;
disk_mem[23466] = 0;
disk_mem[23467] = 0;
disk_mem[23468] = 0;
disk_mem[23469] = 0;
disk_mem[23470] = 0;
disk_mem[23471] = 0;
disk_mem[23472] = 0;
disk_mem[23473] = 0;
disk_mem[23474] = 0;
disk_mem[23475] = 0;
disk_mem[23476] = 0;
disk_mem[23477] = 0;
disk_mem[23478] = 0;
disk_mem[23479] = 0;
disk_mem[23480] = 0;
disk_mem[23481] = 0;
disk_mem[23482] = 0;
disk_mem[23483] = 0;
disk_mem[23484] = 0;
disk_mem[23485] = 0;
disk_mem[23486] = 0;
disk_mem[23487] = 0;
disk_mem[23488] = 0;
disk_mem[23489] = 0;
disk_mem[23490] = 0;
disk_mem[23491] = 0;
disk_mem[23492] = 0;
disk_mem[23493] = 0;
disk_mem[23494] = 0;
disk_mem[23495] = 0;
disk_mem[23496] = 0;
disk_mem[23497] = 0;
disk_mem[23498] = 0;
disk_mem[23499] = 0;
disk_mem[23500] = 0;
disk_mem[23501] = 0;
disk_mem[23502] = 0;
disk_mem[23503] = 0;
disk_mem[23504] = 0;
disk_mem[23505] = 0;
disk_mem[23506] = 0;
disk_mem[23507] = 0;
disk_mem[23508] = 0;
disk_mem[23509] = 0;
disk_mem[23510] = 0;
disk_mem[23511] = 0;
disk_mem[23512] = 0;
disk_mem[23513] = 0;
disk_mem[23514] = 0;
disk_mem[23515] = 0;
disk_mem[23516] = 0;
disk_mem[23517] = 0;
disk_mem[23518] = 0;
disk_mem[23519] = 0;
disk_mem[23520] = 0;
disk_mem[23521] = 0;
disk_mem[23522] = 0;
disk_mem[23523] = 0;
disk_mem[23524] = 0;
disk_mem[23525] = 0;
disk_mem[23526] = 0;
disk_mem[23527] = 0;
disk_mem[23528] = 0;
disk_mem[23529] = 0;
disk_mem[23530] = 0;
disk_mem[23531] = 0;
disk_mem[23532] = 0;
disk_mem[23533] = 0;
disk_mem[23534] = 0;
disk_mem[23535] = 0;
disk_mem[23536] = 0;
disk_mem[23537] = 0;
disk_mem[23538] = 0;
disk_mem[23539] = 0;
disk_mem[23540] = 0;
disk_mem[23541] = 0;
disk_mem[23542] = 0;
disk_mem[23543] = 0;
disk_mem[23544] = 0;
disk_mem[23545] = 0;
disk_mem[23546] = 0;
disk_mem[23547] = 0;
disk_mem[23548] = 0;
disk_mem[23549] = 0;
disk_mem[23550] = 0;
disk_mem[23551] = 0;
disk_mem[23552] = 0;
disk_mem[23553] = 0;
disk_mem[23554] = 0;
disk_mem[23555] = 0;
disk_mem[23556] = 0;
disk_mem[23557] = 0;
disk_mem[23558] = 0;
disk_mem[23559] = 0;
disk_mem[23560] = 0;
disk_mem[23561] = 0;
disk_mem[23562] = 0;
disk_mem[23563] = 0;
disk_mem[23564] = 0;
disk_mem[23565] = 0;
disk_mem[23566] = 0;
disk_mem[23567] = 0;
disk_mem[23568] = 0;
disk_mem[23569] = 0;
disk_mem[23570] = 0;
disk_mem[23571] = 0;
disk_mem[23572] = 0;
disk_mem[23573] = 0;
disk_mem[23574] = 0;
disk_mem[23575] = 0;
disk_mem[23576] = 0;
disk_mem[23577] = 0;
disk_mem[23578] = 0;
disk_mem[23579] = 0;
disk_mem[23580] = 0;
disk_mem[23581] = 0;
disk_mem[23582] = 0;
disk_mem[23583] = 0;
disk_mem[23584] = 0;
disk_mem[23585] = 0;
disk_mem[23586] = 0;
disk_mem[23587] = 0;
disk_mem[23588] = 0;
disk_mem[23589] = 0;
disk_mem[23590] = 0;
disk_mem[23591] = 0;
disk_mem[23592] = 0;
disk_mem[23593] = 0;
disk_mem[23594] = 0;
disk_mem[23595] = 0;
disk_mem[23596] = 0;
disk_mem[23597] = 0;
disk_mem[23598] = 0;
disk_mem[23599] = 0;
disk_mem[23600] = 0;
disk_mem[23601] = 0;
disk_mem[23602] = 0;
disk_mem[23603] = 0;
disk_mem[23604] = 0;
disk_mem[23605] = 0;
disk_mem[23606] = 0;
disk_mem[23607] = 0;
disk_mem[23608] = 0;
disk_mem[23609] = 0;
disk_mem[23610] = 0;
disk_mem[23611] = 0;
disk_mem[23612] = 0;
disk_mem[23613] = 0;
disk_mem[23614] = 0;
disk_mem[23615] = 0;
disk_mem[23616] = 0;
disk_mem[23617] = 0;
disk_mem[23618] = 0;
disk_mem[23619] = 0;
disk_mem[23620] = 0;
disk_mem[23621] = 0;
disk_mem[23622] = 0;
disk_mem[23623] = 0;
disk_mem[23624] = 0;
disk_mem[23625] = 0;
disk_mem[23626] = 0;
disk_mem[23627] = 0;
disk_mem[23628] = 0;
disk_mem[23629] = 0;
disk_mem[23630] = 0;
disk_mem[23631] = 0;
disk_mem[23632] = 0;
disk_mem[23633] = 0;
disk_mem[23634] = 0;
disk_mem[23635] = 0;
disk_mem[23636] = 0;
disk_mem[23637] = 0;
disk_mem[23638] = 0;
disk_mem[23639] = 0;
disk_mem[23640] = 0;
disk_mem[23641] = 0;
disk_mem[23642] = 0;
disk_mem[23643] = 0;
disk_mem[23644] = 0;
disk_mem[23645] = 0;
disk_mem[23646] = 0;
disk_mem[23647] = 0;
disk_mem[23648] = 0;
disk_mem[23649] = 0;
disk_mem[23650] = 0;
disk_mem[23651] = 0;
disk_mem[23652] = 0;
disk_mem[23653] = 0;
disk_mem[23654] = 0;
disk_mem[23655] = 0;
disk_mem[23656] = 0;
disk_mem[23657] = 0;
disk_mem[23658] = 0;
disk_mem[23659] = 0;
disk_mem[23660] = 0;
disk_mem[23661] = 0;
disk_mem[23662] = 0;
disk_mem[23663] = 0;
disk_mem[23664] = 0;
disk_mem[23665] = 0;
disk_mem[23666] = 0;
disk_mem[23667] = 0;
disk_mem[23668] = 0;
disk_mem[23669] = 0;
disk_mem[23670] = 0;
disk_mem[23671] = 0;
disk_mem[23672] = 0;
disk_mem[23673] = 0;
disk_mem[23674] = 0;
disk_mem[23675] = 0;
disk_mem[23676] = 0;
disk_mem[23677] = 0;
disk_mem[23678] = 0;
disk_mem[23679] = 0;
disk_mem[23680] = 0;
disk_mem[23681] = 0;
disk_mem[23682] = 0;
disk_mem[23683] = 0;
disk_mem[23684] = 0;
disk_mem[23685] = 0;
disk_mem[23686] = 0;
disk_mem[23687] = 0;
disk_mem[23688] = 0;
disk_mem[23689] = 0;
disk_mem[23690] = 0;
disk_mem[23691] = 0;
disk_mem[23692] = 0;
disk_mem[23693] = 0;
disk_mem[23694] = 0;
disk_mem[23695] = 0;
disk_mem[23696] = 0;
disk_mem[23697] = 0;
disk_mem[23698] = 0;
disk_mem[23699] = 0;
disk_mem[23700] = 0;
disk_mem[23701] = 0;
disk_mem[23702] = 0;
disk_mem[23703] = 0;
disk_mem[23704] = 0;
disk_mem[23705] = 0;
disk_mem[23706] = 0;
disk_mem[23707] = 0;
disk_mem[23708] = 0;
disk_mem[23709] = 0;
disk_mem[23710] = 0;
disk_mem[23711] = 0;
disk_mem[23712] = 0;
disk_mem[23713] = 0;
disk_mem[23714] = 0;
disk_mem[23715] = 0;
disk_mem[23716] = 0;
disk_mem[23717] = 0;
disk_mem[23718] = 0;
disk_mem[23719] = 0;
disk_mem[23720] = 0;
disk_mem[23721] = 0;
disk_mem[23722] = 0;
disk_mem[23723] = 0;
disk_mem[23724] = 0;
disk_mem[23725] = 0;
disk_mem[23726] = 0;
disk_mem[23727] = 0;
disk_mem[23728] = 0;
disk_mem[23729] = 0;
disk_mem[23730] = 0;
disk_mem[23731] = 0;
disk_mem[23732] = 0;
disk_mem[23733] = 0;
disk_mem[23734] = 0;
disk_mem[23735] = 0;
disk_mem[23736] = 0;
disk_mem[23737] = 0;
disk_mem[23738] = 0;
disk_mem[23739] = 0;
disk_mem[23740] = 0;
disk_mem[23741] = 0;
disk_mem[23742] = 0;
disk_mem[23743] = 0;
disk_mem[23744] = 0;
disk_mem[23745] = 0;
disk_mem[23746] = 0;
disk_mem[23747] = 0;
disk_mem[23748] = 0;
disk_mem[23749] = 0;
disk_mem[23750] = 0;
disk_mem[23751] = 0;
disk_mem[23752] = 0;
disk_mem[23753] = 0;
disk_mem[23754] = 0;
disk_mem[23755] = 0;
disk_mem[23756] = 0;
disk_mem[23757] = 0;
disk_mem[23758] = 0;
disk_mem[23759] = 0;
disk_mem[23760] = 0;
disk_mem[23761] = 0;
disk_mem[23762] = 0;
disk_mem[23763] = 0;
disk_mem[23764] = 0;
disk_mem[23765] = 0;
disk_mem[23766] = 0;
disk_mem[23767] = 0;
disk_mem[23768] = 0;
disk_mem[23769] = 0;
disk_mem[23770] = 0;
disk_mem[23771] = 0;
disk_mem[23772] = 0;
disk_mem[23773] = 0;
disk_mem[23774] = 0;
disk_mem[23775] = 0;
disk_mem[23776] = 0;
disk_mem[23777] = 0;
disk_mem[23778] = 0;
disk_mem[23779] = 0;
disk_mem[23780] = 0;
disk_mem[23781] = 0;
disk_mem[23782] = 0;
disk_mem[23783] = 0;
disk_mem[23784] = 0;
disk_mem[23785] = 0;
disk_mem[23786] = 0;
disk_mem[23787] = 0;
disk_mem[23788] = 0;
disk_mem[23789] = 0;
disk_mem[23790] = 0;
disk_mem[23791] = 0;
disk_mem[23792] = 0;
disk_mem[23793] = 0;
disk_mem[23794] = 0;
disk_mem[23795] = 0;
disk_mem[23796] = 0;
disk_mem[23797] = 0;
disk_mem[23798] = 0;
disk_mem[23799] = 0;
disk_mem[23800] = 0;
disk_mem[23801] = 0;
disk_mem[23802] = 0;
disk_mem[23803] = 0;
disk_mem[23804] = 0;
disk_mem[23805] = 0;
disk_mem[23806] = 0;
disk_mem[23807] = 0;
disk_mem[23808] = 0;
disk_mem[23809] = 0;
disk_mem[23810] = 0;
disk_mem[23811] = 0;
disk_mem[23812] = 0;
disk_mem[23813] = 0;
disk_mem[23814] = 0;
disk_mem[23815] = 0;
disk_mem[23816] = 0;
disk_mem[23817] = 0;
disk_mem[23818] = 0;
disk_mem[23819] = 0;
disk_mem[23820] = 0;
disk_mem[23821] = 0;
disk_mem[23822] = 0;
disk_mem[23823] = 0;
disk_mem[23824] = 0;
disk_mem[23825] = 0;
disk_mem[23826] = 0;
disk_mem[23827] = 0;
disk_mem[23828] = 0;
disk_mem[23829] = 0;
disk_mem[23830] = 0;
disk_mem[23831] = 0;
disk_mem[23832] = 0;
disk_mem[23833] = 0;
disk_mem[23834] = 0;
disk_mem[23835] = 0;
disk_mem[23836] = 0;
disk_mem[23837] = 0;
disk_mem[23838] = 0;
disk_mem[23839] = 0;
disk_mem[23840] = 0;
disk_mem[23841] = 0;
disk_mem[23842] = 0;
disk_mem[23843] = 0;
disk_mem[23844] = 0;
disk_mem[23845] = 0;
disk_mem[23846] = 0;
disk_mem[23847] = 0;
disk_mem[23848] = 0;
disk_mem[23849] = 0;
disk_mem[23850] = 0;
disk_mem[23851] = 0;
disk_mem[23852] = 0;
disk_mem[23853] = 0;
disk_mem[23854] = 0;
disk_mem[23855] = 0;
disk_mem[23856] = 0;
disk_mem[23857] = 0;
disk_mem[23858] = 0;
disk_mem[23859] = 0;
disk_mem[23860] = 0;
disk_mem[23861] = 0;
disk_mem[23862] = 0;
disk_mem[23863] = 0;
disk_mem[23864] = 0;
disk_mem[23865] = 0;
disk_mem[23866] = 0;
disk_mem[23867] = 0;
disk_mem[23868] = 0;
disk_mem[23869] = 0;
disk_mem[23870] = 0;
disk_mem[23871] = 0;
disk_mem[23872] = 0;
disk_mem[23873] = 0;
disk_mem[23874] = 0;
disk_mem[23875] = 0;
disk_mem[23876] = 0;
disk_mem[23877] = 0;
disk_mem[23878] = 0;
disk_mem[23879] = 0;
disk_mem[23880] = 0;
disk_mem[23881] = 0;
disk_mem[23882] = 0;
disk_mem[23883] = 0;
disk_mem[23884] = 0;
disk_mem[23885] = 0;
disk_mem[23886] = 0;
disk_mem[23887] = 0;
disk_mem[23888] = 0;
disk_mem[23889] = 0;
disk_mem[23890] = 0;
disk_mem[23891] = 0;
disk_mem[23892] = 0;
disk_mem[23893] = 0;
disk_mem[23894] = 0;
disk_mem[23895] = 0;
disk_mem[23896] = 0;
disk_mem[23897] = 0;
disk_mem[23898] = 0;
disk_mem[23899] = 0;
disk_mem[23900] = 0;
disk_mem[23901] = 0;
disk_mem[23902] = 0;
disk_mem[23903] = 0;
disk_mem[23904] = 0;
disk_mem[23905] = 0;
disk_mem[23906] = 0;
disk_mem[23907] = 0;
disk_mem[23908] = 0;
disk_mem[23909] = 0;
disk_mem[23910] = 0;
disk_mem[23911] = 0;
disk_mem[23912] = 0;
disk_mem[23913] = 0;
disk_mem[23914] = 0;
disk_mem[23915] = 0;
disk_mem[23916] = 0;
disk_mem[23917] = 0;
disk_mem[23918] = 0;
disk_mem[23919] = 0;
disk_mem[23920] = 0;
disk_mem[23921] = 0;
disk_mem[23922] = 0;
disk_mem[23923] = 0;
disk_mem[23924] = 0;
disk_mem[23925] = 0;
disk_mem[23926] = 0;
disk_mem[23927] = 0;
disk_mem[23928] = 0;
disk_mem[23929] = 0;
disk_mem[23930] = 0;
disk_mem[23931] = 0;
disk_mem[23932] = 0;
disk_mem[23933] = 0;
disk_mem[23934] = 0;
disk_mem[23935] = 0;
disk_mem[23936] = 0;
disk_mem[23937] = 0;
disk_mem[23938] = 0;
disk_mem[23939] = 0;
disk_mem[23940] = 0;
disk_mem[23941] = 0;
disk_mem[23942] = 0;
disk_mem[23943] = 0;
disk_mem[23944] = 0;
disk_mem[23945] = 0;
disk_mem[23946] = 0;
disk_mem[23947] = 0;
disk_mem[23948] = 0;
disk_mem[23949] = 0;
disk_mem[23950] = 0;
disk_mem[23951] = 0;
disk_mem[23952] = 0;
disk_mem[23953] = 0;
disk_mem[23954] = 0;
disk_mem[23955] = 0;
disk_mem[23956] = 0;
disk_mem[23957] = 0;
disk_mem[23958] = 0;
disk_mem[23959] = 0;
disk_mem[23960] = 0;
disk_mem[23961] = 0;
disk_mem[23962] = 0;
disk_mem[23963] = 0;
disk_mem[23964] = 0;
disk_mem[23965] = 0;
disk_mem[23966] = 0;
disk_mem[23967] = 0;
disk_mem[23968] = 0;
disk_mem[23969] = 0;
disk_mem[23970] = 0;
disk_mem[23971] = 0;
disk_mem[23972] = 0;
disk_mem[23973] = 0;
disk_mem[23974] = 0;
disk_mem[23975] = 0;
disk_mem[23976] = 0;
disk_mem[23977] = 0;
disk_mem[23978] = 0;
disk_mem[23979] = 0;
disk_mem[23980] = 0;
disk_mem[23981] = 0;
disk_mem[23982] = 0;
disk_mem[23983] = 0;
disk_mem[23984] = 0;
disk_mem[23985] = 0;
disk_mem[23986] = 0;
disk_mem[23987] = 0;
disk_mem[23988] = 0;
disk_mem[23989] = 0;
disk_mem[23990] = 0;
disk_mem[23991] = 0;
disk_mem[23992] = 0;
disk_mem[23993] = 0;
disk_mem[23994] = 0;
disk_mem[23995] = 0;
disk_mem[23996] = 0;
disk_mem[23997] = 0;
disk_mem[23998] = 0;
disk_mem[23999] = 0;
disk_mem[24000] = 0;
disk_mem[24001] = 0;
disk_mem[24002] = 0;
disk_mem[24003] = 0;
disk_mem[24004] = 0;
disk_mem[24005] = 0;
disk_mem[24006] = 0;
disk_mem[24007] = 0;
disk_mem[24008] = 0;
disk_mem[24009] = 0;
disk_mem[24010] = 0;
disk_mem[24011] = 0;
disk_mem[24012] = 0;
disk_mem[24013] = 0;
disk_mem[24014] = 0;
disk_mem[24015] = 0;
disk_mem[24016] = 0;
disk_mem[24017] = 0;
disk_mem[24018] = 0;
disk_mem[24019] = 0;
disk_mem[24020] = 0;
disk_mem[24021] = 0;
disk_mem[24022] = 0;
disk_mem[24023] = 0;
disk_mem[24024] = 0;
disk_mem[24025] = 0;
disk_mem[24026] = 0;
disk_mem[24027] = 0;
disk_mem[24028] = 0;
disk_mem[24029] = 0;
disk_mem[24030] = 0;
disk_mem[24031] = 0;
disk_mem[24032] = 0;
disk_mem[24033] = 0;
disk_mem[24034] = 0;
disk_mem[24035] = 0;
disk_mem[24036] = 0;
disk_mem[24037] = 0;
disk_mem[24038] = 0;
disk_mem[24039] = 0;
disk_mem[24040] = 0;
disk_mem[24041] = 0;
disk_mem[24042] = 0;
disk_mem[24043] = 0;
disk_mem[24044] = 0;
disk_mem[24045] = 0;
disk_mem[24046] = 0;
disk_mem[24047] = 0;
disk_mem[24048] = 0;
disk_mem[24049] = 0;
disk_mem[24050] = 0;
disk_mem[24051] = 0;
disk_mem[24052] = 0;
disk_mem[24053] = 0;
disk_mem[24054] = 0;
disk_mem[24055] = 0;
disk_mem[24056] = 0;
disk_mem[24057] = 0;
disk_mem[24058] = 0;
disk_mem[24059] = 0;
disk_mem[24060] = 0;
disk_mem[24061] = 0;
disk_mem[24062] = 0;
disk_mem[24063] = 0;
disk_mem[24064] = 0;
disk_mem[24065] = 0;
disk_mem[24066] = 0;
disk_mem[24067] = 0;
disk_mem[24068] = 0;
disk_mem[24069] = 0;
disk_mem[24070] = 0;
disk_mem[24071] = 0;
disk_mem[24072] = 0;
disk_mem[24073] = 0;
disk_mem[24074] = 0;
disk_mem[24075] = 0;
disk_mem[24076] = 0;
disk_mem[24077] = 0;
disk_mem[24078] = 0;
disk_mem[24079] = 0;
disk_mem[24080] = 0;
disk_mem[24081] = 0;
disk_mem[24082] = 0;
disk_mem[24083] = 0;
disk_mem[24084] = 0;
disk_mem[24085] = 0;
disk_mem[24086] = 0;
disk_mem[24087] = 0;
disk_mem[24088] = 0;
disk_mem[24089] = 0;
disk_mem[24090] = 0;
disk_mem[24091] = 0;
disk_mem[24092] = 0;
disk_mem[24093] = 0;
disk_mem[24094] = 0;
disk_mem[24095] = 0;
disk_mem[24096] = 0;
disk_mem[24097] = 0;
disk_mem[24098] = 0;
disk_mem[24099] = 0;
disk_mem[24100] = 0;
disk_mem[24101] = 0;
disk_mem[24102] = 0;
disk_mem[24103] = 0;
disk_mem[24104] = 0;
disk_mem[24105] = 0;
disk_mem[24106] = 0;
disk_mem[24107] = 0;
disk_mem[24108] = 0;
disk_mem[24109] = 0;
disk_mem[24110] = 0;
disk_mem[24111] = 0;
disk_mem[24112] = 0;
disk_mem[24113] = 0;
disk_mem[24114] = 0;
disk_mem[24115] = 0;
disk_mem[24116] = 0;
disk_mem[24117] = 0;
disk_mem[24118] = 0;
disk_mem[24119] = 0;
disk_mem[24120] = 0;
disk_mem[24121] = 0;
disk_mem[24122] = 0;
disk_mem[24123] = 0;
disk_mem[24124] = 0;
disk_mem[24125] = 0;
disk_mem[24126] = 0;
disk_mem[24127] = 0;
disk_mem[24128] = 0;
disk_mem[24129] = 0;
disk_mem[24130] = 0;
disk_mem[24131] = 0;
disk_mem[24132] = 0;
disk_mem[24133] = 0;
disk_mem[24134] = 0;
disk_mem[24135] = 0;
disk_mem[24136] = 0;
disk_mem[24137] = 0;
disk_mem[24138] = 0;
disk_mem[24139] = 0;
disk_mem[24140] = 0;
disk_mem[24141] = 0;
disk_mem[24142] = 0;
disk_mem[24143] = 0;
disk_mem[24144] = 0;
disk_mem[24145] = 0;
disk_mem[24146] = 0;
disk_mem[24147] = 0;
disk_mem[24148] = 0;
disk_mem[24149] = 0;
disk_mem[24150] = 0;
disk_mem[24151] = 0;
disk_mem[24152] = 0;
disk_mem[24153] = 0;
disk_mem[24154] = 0;
disk_mem[24155] = 0;
disk_mem[24156] = 0;
disk_mem[24157] = 0;
disk_mem[24158] = 0;
disk_mem[24159] = 0;
disk_mem[24160] = 0;
disk_mem[24161] = 0;
disk_mem[24162] = 0;
disk_mem[24163] = 0;
disk_mem[24164] = 0;
disk_mem[24165] = 0;
disk_mem[24166] = 0;
disk_mem[24167] = 0;
disk_mem[24168] = 0;
disk_mem[24169] = 0;
disk_mem[24170] = 0;
disk_mem[24171] = 0;
disk_mem[24172] = 0;
disk_mem[24173] = 0;
disk_mem[24174] = 0;
disk_mem[24175] = 0;
disk_mem[24176] = 0;
disk_mem[24177] = 0;
disk_mem[24178] = 0;
disk_mem[24179] = 0;
disk_mem[24180] = 0;
disk_mem[24181] = 0;
disk_mem[24182] = 0;
disk_mem[24183] = 0;
disk_mem[24184] = 0;
disk_mem[24185] = 0;
disk_mem[24186] = 0;
disk_mem[24187] = 0;
disk_mem[24188] = 0;
disk_mem[24189] = 0;
disk_mem[24190] = 0;
disk_mem[24191] = 0;
disk_mem[24192] = 0;
disk_mem[24193] = 0;
disk_mem[24194] = 0;
disk_mem[24195] = 0;
disk_mem[24196] = 0;
disk_mem[24197] = 0;
disk_mem[24198] = 0;
disk_mem[24199] = 0;
disk_mem[24200] = 0;
disk_mem[24201] = 0;
disk_mem[24202] = 0;
disk_mem[24203] = 0;
disk_mem[24204] = 0;
disk_mem[24205] = 0;
disk_mem[24206] = 0;
disk_mem[24207] = 0;
disk_mem[24208] = 0;
disk_mem[24209] = 0;
disk_mem[24210] = 0;
disk_mem[24211] = 0;
disk_mem[24212] = 0;
disk_mem[24213] = 0;
disk_mem[24214] = 0;
disk_mem[24215] = 0;
disk_mem[24216] = 0;
disk_mem[24217] = 0;
disk_mem[24218] = 0;
disk_mem[24219] = 0;
disk_mem[24220] = 0;
disk_mem[24221] = 0;
disk_mem[24222] = 0;
disk_mem[24223] = 0;
disk_mem[24224] = 0;
disk_mem[24225] = 0;
disk_mem[24226] = 0;
disk_mem[24227] = 0;
disk_mem[24228] = 0;
disk_mem[24229] = 0;
disk_mem[24230] = 0;
disk_mem[24231] = 0;
disk_mem[24232] = 0;
disk_mem[24233] = 0;
disk_mem[24234] = 0;
disk_mem[24235] = 0;
disk_mem[24236] = 0;
disk_mem[24237] = 0;
disk_mem[24238] = 0;
disk_mem[24239] = 0;
disk_mem[24240] = 0;
disk_mem[24241] = 0;
disk_mem[24242] = 0;
disk_mem[24243] = 0;
disk_mem[24244] = 0;
disk_mem[24245] = 0;
disk_mem[24246] = 0;
disk_mem[24247] = 0;
disk_mem[24248] = 0;
disk_mem[24249] = 0;
disk_mem[24250] = 0;
disk_mem[24251] = 0;
disk_mem[24252] = 0;
disk_mem[24253] = 0;
disk_mem[24254] = 0;
disk_mem[24255] = 0;
disk_mem[24256] = 0;
disk_mem[24257] = 0;
disk_mem[24258] = 0;
disk_mem[24259] = 0;
disk_mem[24260] = 0;
disk_mem[24261] = 0;
disk_mem[24262] = 0;
disk_mem[24263] = 0;
disk_mem[24264] = 0;
disk_mem[24265] = 0;
disk_mem[24266] = 0;
disk_mem[24267] = 0;
disk_mem[24268] = 0;
disk_mem[24269] = 0;
disk_mem[24270] = 0;
disk_mem[24271] = 0;
disk_mem[24272] = 0;
disk_mem[24273] = 0;
disk_mem[24274] = 0;
disk_mem[24275] = 0;
disk_mem[24276] = 0;
disk_mem[24277] = 0;
disk_mem[24278] = 0;
disk_mem[24279] = 0;
disk_mem[24280] = 0;
disk_mem[24281] = 0;
disk_mem[24282] = 0;
disk_mem[24283] = 0;
disk_mem[24284] = 0;
disk_mem[24285] = 0;
disk_mem[24286] = 0;
disk_mem[24287] = 0;
disk_mem[24288] = 0;
disk_mem[24289] = 0;
disk_mem[24290] = 0;
disk_mem[24291] = 0;
disk_mem[24292] = 0;
disk_mem[24293] = 0;
disk_mem[24294] = 0;
disk_mem[24295] = 0;
disk_mem[24296] = 0;
disk_mem[24297] = 0;
disk_mem[24298] = 0;
disk_mem[24299] = 0;
disk_mem[24300] = 0;
disk_mem[24301] = 0;
disk_mem[24302] = 0;
disk_mem[24303] = 0;
disk_mem[24304] = 0;
disk_mem[24305] = 0;
disk_mem[24306] = 0;
disk_mem[24307] = 0;
disk_mem[24308] = 0;
disk_mem[24309] = 0;
disk_mem[24310] = 0;
disk_mem[24311] = 0;
disk_mem[24312] = 0;
disk_mem[24313] = 0;
disk_mem[24314] = 0;
disk_mem[24315] = 0;
disk_mem[24316] = 0;
disk_mem[24317] = 0;
disk_mem[24318] = 0;
disk_mem[24319] = 0;
disk_mem[24320] = 0;
disk_mem[24321] = 0;
disk_mem[24322] = 0;
disk_mem[24323] = 0;
disk_mem[24324] = 0;
disk_mem[24325] = 0;
disk_mem[24326] = 0;
disk_mem[24327] = 0;
disk_mem[24328] = 0;
disk_mem[24329] = 0;
disk_mem[24330] = 0;
disk_mem[24331] = 0;
disk_mem[24332] = 0;
disk_mem[24333] = 0;
disk_mem[24334] = 0;
disk_mem[24335] = 0;
disk_mem[24336] = 0;
disk_mem[24337] = 0;
disk_mem[24338] = 0;
disk_mem[24339] = 0;
disk_mem[24340] = 0;
disk_mem[24341] = 0;
disk_mem[24342] = 0;
disk_mem[24343] = 0;
disk_mem[24344] = 0;
disk_mem[24345] = 0;
disk_mem[24346] = 0;
disk_mem[24347] = 0;
disk_mem[24348] = 0;
disk_mem[24349] = 0;
disk_mem[24350] = 0;
disk_mem[24351] = 0;
disk_mem[24352] = 0;
disk_mem[24353] = 0;
disk_mem[24354] = 0;
disk_mem[24355] = 0;
disk_mem[24356] = 0;
disk_mem[24357] = 0;
disk_mem[24358] = 0;
disk_mem[24359] = 0;
disk_mem[24360] = 0;
disk_mem[24361] = 0;
disk_mem[24362] = 0;
disk_mem[24363] = 0;
disk_mem[24364] = 0;
disk_mem[24365] = 0;
disk_mem[24366] = 0;
disk_mem[24367] = 0;
disk_mem[24368] = 0;
disk_mem[24369] = 0;
disk_mem[24370] = 0;
disk_mem[24371] = 0;
disk_mem[24372] = 0;
disk_mem[24373] = 0;
disk_mem[24374] = 0;
disk_mem[24375] = 0;
disk_mem[24376] = 0;
disk_mem[24377] = 0;
disk_mem[24378] = 0;
disk_mem[24379] = 0;
disk_mem[24380] = 0;
disk_mem[24381] = 0;
disk_mem[24382] = 0;
disk_mem[24383] = 0;
disk_mem[24384] = 0;
disk_mem[24385] = 0;
disk_mem[24386] = 0;
disk_mem[24387] = 0;
disk_mem[24388] = 0;
disk_mem[24389] = 0;
disk_mem[24390] = 0;
disk_mem[24391] = 0;
disk_mem[24392] = 0;
disk_mem[24393] = 0;
disk_mem[24394] = 0;
disk_mem[24395] = 0;
disk_mem[24396] = 0;
disk_mem[24397] = 0;
disk_mem[24398] = 0;
disk_mem[24399] = 0;
disk_mem[24400] = 0;
disk_mem[24401] = 0;
disk_mem[24402] = 0;
disk_mem[24403] = 0;
disk_mem[24404] = 0;
disk_mem[24405] = 0;
disk_mem[24406] = 0;
disk_mem[24407] = 0;
disk_mem[24408] = 0;
disk_mem[24409] = 0;
disk_mem[24410] = 0;
disk_mem[24411] = 0;
disk_mem[24412] = 0;
disk_mem[24413] = 0;
disk_mem[24414] = 0;
disk_mem[24415] = 0;
disk_mem[24416] = 0;
disk_mem[24417] = 0;
disk_mem[24418] = 0;
disk_mem[24419] = 0;
disk_mem[24420] = 0;
disk_mem[24421] = 0;
disk_mem[24422] = 0;
disk_mem[24423] = 0;
disk_mem[24424] = 0;
disk_mem[24425] = 0;
disk_mem[24426] = 0;
disk_mem[24427] = 0;
disk_mem[24428] = 0;
disk_mem[24429] = 0;
disk_mem[24430] = 0;
disk_mem[24431] = 0;
disk_mem[24432] = 0;
disk_mem[24433] = 0;
disk_mem[24434] = 0;
disk_mem[24435] = 0;
disk_mem[24436] = 0;
disk_mem[24437] = 0;
disk_mem[24438] = 0;
disk_mem[24439] = 0;
disk_mem[24440] = 0;
disk_mem[24441] = 0;
disk_mem[24442] = 0;
disk_mem[24443] = 0;
disk_mem[24444] = 0;
disk_mem[24445] = 0;
disk_mem[24446] = 0;
disk_mem[24447] = 0;
disk_mem[24448] = 0;
disk_mem[24449] = 0;
disk_mem[24450] = 0;
disk_mem[24451] = 0;
disk_mem[24452] = 0;
disk_mem[24453] = 0;
disk_mem[24454] = 0;
disk_mem[24455] = 0;
disk_mem[24456] = 0;
disk_mem[24457] = 0;
disk_mem[24458] = 0;
disk_mem[24459] = 0;
disk_mem[24460] = 0;
disk_mem[24461] = 0;
disk_mem[24462] = 0;
disk_mem[24463] = 0;
disk_mem[24464] = 0;
disk_mem[24465] = 0;
disk_mem[24466] = 0;
disk_mem[24467] = 0;
disk_mem[24468] = 0;
disk_mem[24469] = 0;
disk_mem[24470] = 0;
disk_mem[24471] = 0;
disk_mem[24472] = 0;
disk_mem[24473] = 0;
disk_mem[24474] = 0;
disk_mem[24475] = 0;
disk_mem[24476] = 0;
disk_mem[24477] = 0;
disk_mem[24478] = 0;
disk_mem[24479] = 0;
disk_mem[24480] = 0;
disk_mem[24481] = 0;
disk_mem[24482] = 0;
disk_mem[24483] = 0;
disk_mem[24484] = 0;
disk_mem[24485] = 0;
disk_mem[24486] = 0;
disk_mem[24487] = 0;
disk_mem[24488] = 0;
disk_mem[24489] = 0;
disk_mem[24490] = 0;
disk_mem[24491] = 0;
disk_mem[24492] = 0;
disk_mem[24493] = 0;
disk_mem[24494] = 0;
disk_mem[24495] = 0;
disk_mem[24496] = 0;
disk_mem[24497] = 0;
disk_mem[24498] = 0;
disk_mem[24499] = 0;
disk_mem[24500] = 0;
disk_mem[24501] = 0;
disk_mem[24502] = 0;
disk_mem[24503] = 0;
disk_mem[24504] = 0;
disk_mem[24505] = 0;
disk_mem[24506] = 0;
disk_mem[24507] = 0;
disk_mem[24508] = 0;
disk_mem[24509] = 0;
disk_mem[24510] = 0;
disk_mem[24511] = 0;
disk_mem[24512] = 0;
disk_mem[24513] = 0;
disk_mem[24514] = 0;
disk_mem[24515] = 0;
disk_mem[24516] = 0;
disk_mem[24517] = 0;
disk_mem[24518] = 0;
disk_mem[24519] = 0;
disk_mem[24520] = 0;
disk_mem[24521] = 0;
disk_mem[24522] = 0;
disk_mem[24523] = 0;
disk_mem[24524] = 0;
disk_mem[24525] = 0;
disk_mem[24526] = 0;
disk_mem[24527] = 0;
disk_mem[24528] = 0;
disk_mem[24529] = 0;
disk_mem[24530] = 0;
disk_mem[24531] = 0;
disk_mem[24532] = 0;
disk_mem[24533] = 0;
disk_mem[24534] = 0;
disk_mem[24535] = 0;
disk_mem[24536] = 0;
disk_mem[24537] = 0;
disk_mem[24538] = 0;
disk_mem[24539] = 0;
disk_mem[24540] = 0;
disk_mem[24541] = 0;
disk_mem[24542] = 0;
disk_mem[24543] = 0;
disk_mem[24544] = 0;
disk_mem[24545] = 0;
disk_mem[24546] = 0;
disk_mem[24547] = 0;
disk_mem[24548] = 0;
disk_mem[24549] = 0;
disk_mem[24550] = 0;
disk_mem[24551] = 0;
disk_mem[24552] = 0;
disk_mem[24553] = 0;
disk_mem[24554] = 0;
disk_mem[24555] = 0;
disk_mem[24556] = 0;
disk_mem[24557] = 0;
disk_mem[24558] = 0;
disk_mem[24559] = 0;
disk_mem[24560] = 0;
disk_mem[24561] = 0;
disk_mem[24562] = 0;
disk_mem[24563] = 0;
disk_mem[24564] = 0;
disk_mem[24565] = 0;
disk_mem[24566] = 0;
disk_mem[24567] = 0;
disk_mem[24568] = 0;
disk_mem[24569] = 0;
disk_mem[24570] = 0;
disk_mem[24571] = 0;
disk_mem[24572] = 0;
disk_mem[24573] = 0;
disk_mem[24574] = 0;
disk_mem[24575] = 0;
end


endmodule
